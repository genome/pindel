#COLO-829_BL.bam	mean:197.060	std:21.090	uppercutoff:282.340	lowercutoff:113.570	readlen:75.000	library:COLO-829BL-IL	reflen:62427936	seqcov:37.923x	phycov:49.821x	1:756	2:6732	3:36330	4:5916	8:806	32:43397
#COLO-829.bam	mean:456.450	std:22.420	uppercutoff:531.160	lowercutoff:350.560	readlen:36.290	library:COLO-829_v2_74	reflen:62427936	seqcov:2.837x	phycov:17.843x	1:390	2:2904	3:136706	4:1022	8:362	32:32168
#COLO-829.bam	mean:203.220	std:21.370	uppercutoff:287.940	lowercutoff:116.960	readlen:75.000	library:COLO-829-IL	reflen:62427936	seqcov:60.325x	phycov:81.728x	1:2590	2:11482	3:58012	4:11448	8:2420	32:91908
#Chr1	Pos1	Orientation1	Chr2	Pos2	Orientation2	Type	Size	Score	num_Reads	num_Reads_lib	Allele_frequency	Version	Run_Param
20	21285	2+2-	20	21246	2+2-	INS	-110	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39618	3+3-	20	39670	3+3-	INS	-278	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43162	3+2-	20	43154	3+2-	INS	-94	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47475	2+2-	20	47445	2+2-	INS	-110	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51541	2+2-	20	51585	2+2-	INS	-386	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57076	2+2-	20	57126	2+2-	INS	-104	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	64915	4+2-	20	64976	4+2-	INS	-93	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	69639	2+0-	20	69759	0+2-	INS	-200	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	109762	2+3-	20	109782	2+3-	INS	-104	29	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	111723	2+3-	20	111741	2+3-	INS	-103	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	123027	3+4-	20	123070	3+4-	INS	-194	29	3	COLO-829_v2_74|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	134019	2+2-	20	133989	2+2-	INS	-98	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	134164	2+2-	20	134186	2+2-	INS	-97	28	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	136149	2+1-	20	136196	0+2-	INS	-273	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	136736	2+1-	20	136809	1+4-	INS	-182	30	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	142982	3+0-	20	145331	1+2-	DEL	2306	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	173578	4+3-	20	173580	4+3-	INS	-272	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	174374	3+2-	20	174359	3+2-	INS	-387	21	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	193011	2+2-	20	193030	2+2-	INS	-89	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	214666	4+2-	20	214676	4+2-	INS	-234	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	214746	2+0-	20	214831	1+2-	INS	-223	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	234783	3+0-	20	234901	17+22-	INS	-160	33	6	COLO-829_v2_74|5:COLO-829-IL|1	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	234885	2+0-	20	234901	10+12-	INS	-228	7	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	245847	3+4-	20	245866	3+4-	INS	-103	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	264807	4+6-	20	264861	4+6-	INS	-101	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	278057	2+0-	20	278099	0+2-	INS	-283	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	293666	2+2-	20	293635	2+2-	INS	-119	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	305586	5+3-	20	305591	2+3-	INS	-167	33	5	COLO-829_v2_74|2:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	312429	3+3-	20	312423	3+3-	INS	-272	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	330235	3+0-	20	330363	2+5-	INS	-145	36	4	COLO-829BL-IL|2:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	338030	3+0-	20	338034	0+3-	INS	-299	32	3	COLO-829_v2_74|3	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	373114	2+2-	20	373058	2+2-	INS	-406	33	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	386515	3+2-	20	386534	3+2-	INS	-102	29	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	396718	3+3-	20	396749	3+3-	INS	-100	36	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	399186	11+0-	20	399257	0+16-	INS	-272	12	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	421196	2+2-	20	421157	2+2-	INS	-124	33	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	423563	2+2-	20	423565	2+2-	INS	-94	30	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	435500	2+2-	20	435518	2+2-	INS	-102	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	443070	3+3-	20	443086	3+3-	INS	-102	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	463337	4+3-	20	463396	4+3-	INS	-97	36	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	491154	2+2-	20	491173	2+2-	INS	-94	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	514313	2+3-	20	514353	2+3-	INS	-247	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	514750	2+6-	20	514800	2+6-	INS	-105	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	553215	2+2-	20	553245	2+2-	INS	-394	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	561311	2+0-	20	561497	0+2-	INS	-135	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	577611	2+3-	20	577646	2+3-	INS	-368	16	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	579426	3+2-	20	579395	3+2-	INS	-123	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	588703	2+0-	20	588796	1+2-	INS	-232	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	596353	3+3-	20	596391	3+3-	INS	-171	33	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	600647	2+2-	20	600617	2+2-	INS	-253	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	628017	3+4-	20	628007	3+4-	INS	-107	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	638468	14+0-	20	638522	0+14-	DEL	99	99	12	COLO-829BL-IL|6:COLO-829-IL|6	0.31	BreakDancerMax-0.0.1r81	|q10|o20
20	666799	4+3-	20	666807	4+3-	INS	-253	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	669118	2+0-	20	669179	0+2-	INS	-251	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	669735	4+4-	20	669812	4+4-	INS	-107	20	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	686680	2+2-	20	686634	2+2-	INS	-395	28	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	712851	7+2-	20	712894	7+2-	INS	-101	23	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	718134	2+3-	20	718212	2+3-	INS	-102	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	725225	3+2-	20	725184	3+2-	INS	-109	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	732063	2+3-	20	732034	2+3-	INS	-104	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	767199	2+2-	20	767202	2+2-	INS	-109	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	771303	4+5-	20	771405	4+5-	INS	-105	42	4	COLO-829BL-IL|1:COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	786385	2+2-	20	786352	2+2-	INS	-116	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	787428	3+2-	20	787452	3+2-	INS	-94	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	791363	2+2-	20	791357	2+2-	INS	-100	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	799585	2+0-	20	799671	0+3-	INS	-228	19	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	832888	2+4-	20	832897	2+4-	INS	-90	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	838664	4+2-	20	838703	4+2-	INS	-105	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	838773	2+0-	20	838928	2+4-	INS	-136	27	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	865384	2+0-	20	865442	0+2-	INS	-256	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	878220	19+0-	20	878294	0+21-	DEL	100	99	19	COLO-829BL-IL|9:COLO-829-IL|10	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	886833	2+2-	20	886840	2+2-	INS	-108	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	910443	2+2-	20	910435	2+2-	INS	-98	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	913645	5+2-	20	913707	11+8-	ITX	-138	99	6	COLO-829BL-IL|3:COLO-829-IL|3	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	913645	3+1-	20	913964	0+6-	DEL	277	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	913830	4+0-	20	913964	0+4-	DEL	149	77	4	COLO-829BL-IL|2:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	917413	2+3-	20	917433	2+3-	INS	-98	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	923281	3+3-	20	923317	3+3-	INS	-230	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	927905	2+0-	20	927939	0+2-	INS	-284	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	937726	2+2-	20	937726	2+2-	INS	-92	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	948364	2+0-	20	948494	1+3-	DEL	111	34	2	COLO-829-IL|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	959517	2+2-	20	959535	2+2-	INS	-210	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	989903	2+2-	20	989858	2+2-	INS	-112	35	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1001123	2+2-	20	1001070	2+2-	INS	-402	31	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1016422	2+2-	20	1016415	2+2-	INS	-251	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1021121	2+3-	20	1021115	2+3-	INS	-114	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1023013	2+2-	20	1022992	2+2-	INS	-248	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1028659	13+2-	20	1028735	13+2-	INS	-101	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	1045733	2+2-	20	1045754	2+2-	INS	-103	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1048679	2+2-	20	1048645	2+2-	INS	-255	27	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1055563	2+2-	20	1055553	2+2-	INS	-102	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1060887	3+0-	20	1060911	1+4-	INS	-281	27	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	1069496	4+1-	20	1069533	0+3-	INS	-209	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1072151	3+1-	20	1072216	3+4-	INS	-159	45	5	COLO-829BL-IL|2:COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	1077932	2+3-	20	1077942	2+3-	INS	-231	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1078533	6+3-	20	1078534	6+3-	INS	-120	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1078604	3+0-	20	1078787	2+4-	DEL	92	53	3	COLO-829-IL|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	1087378	2+0-	20	1087434	1+2-	INS	-270	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1095359	2+2-	20	1095312	2+2-	INS	-397	29	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1097867	2+0-	20	1098009	0+2-	INS	-172	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1106226	2+2-	20	1106225	2+2-	INS	-104	27	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1111815	3+3-	20	1111838	3+3-	INS	-99	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1122745	2+3-	20	1122779	2+3-	INS	-204	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1124545	2+2-	20	1124572	2+2-	INS	-93	28	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1133281	2+3-	20	1133261	2+3-	INS	-267	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1138279	3+1-	20	1138355	1+2-	INS	-167	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1158911	3+2-	20	1158933	0+2-	INS	-235	23	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1167912	2+2-	20	1167862	2+2-	INS	-117	37	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1182576	2+4-	20	1182566	2+4-	INS	-111	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1183096	2+3-	20	1183088	2+3-	INS	-97	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1185551	2+2-	20	1185491	2+2-	INS	-121	43	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1189762	2+2-	20	1189753	2+2-	INS	-106	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1197232	2+2-	20	1197216	2+2-	INS	-121	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1206273	2+2-	20	1206256	2+2-	ITX	-178	43	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1210822	2+2-	20	1210824	2+2-	INS	-97	30	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1220522	2+3-	20	1220534	2+3-	INS	-99	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1221429	2+2-	20	1221452	2+2-	INS	-236	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1225947	2+0-	20	1226121	0+2-	INS	-139	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1284077	2+2-	20	1284132	2+2-	INS	-360	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1300207	2+0-	20	1300258	1+4-	INS	-131	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1309053	5+6-	20	1309182	5+6-	INS	-171	31	4	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1327346	6+2-	20	1327415	6+2-	INS	-253	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1328930	2+2-	20	1328945	2+2-	INS	-252	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1336845	3+2-	20	1338811	1+18-	INS	-99	23	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1337164	20+0-	20	1338811	0+15-	DEL	1680	99	15	COLO-829BL-IL|7:COLO-829-IL|8	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	1337164	5+0-	20	1339093	1+5-	DEL	1668	93	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1345617	3+3-	20	1345645	3+3-	INS	-103	38	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1350934	2+2-	20	1350899	2+2-	INS	-385	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1358904	2+2-	20	1358861	2+2-	INS	-100	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1361467	3+2-	20	1361627	1+3-	INS	-152	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1361878	4+4-	20	1362003	4+4-	INS	-354	11	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1399933	3+2-	20	1399958	3+2-	INS	-97	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1403120	5+2-	20	1403169	5+2-	INS	-103	26	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1413739	2+2-	20	1413700	2+2-	INS	-105	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	1414150	2+2-	20	1414153	2+2-	INS	-106	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1439727	3+3-	20	1439760	3+3-	INS	-104	35	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1453748	2+4-	20	1453796	2+4-	INS	-100	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1460947	2+3-	20	1460926	2+3-	INS	-371	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1463326	2+3-	20	1463337	2+3-	INS	-110	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1467005	3+5-	20	1467013	3+5-	INS	-361	31	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1469538	2+2-	20	1469530	2+2-	INS	-107	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1481165	2+2-	20	1481170	2+2-	INS	-112	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1482075	2+2-	20	1482117	2+2-	INS	-226	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1484229	2+2-	20	1484295	2+2-	INS	-92	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1486234	2+2-	20	1486215	2+2-	INS	-100	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1508971	3+1-	20	1542301	0+3-	DEL	33060	48	2	COLO-829_v2_74|2	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	1533438	0+5-	20	1564658	5+0-	ITX	31040	99	5	COLO-829BL-IL|3:COLO-829-IL|2	0.50	BreakDancerMax-0.0.1r81	|q10|o20
20	1550220	2+4-	20	1550306	2+4-	INS	-111	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1551237	2+2-	20	1551227	2+2-	INS	-105	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1596864	12+4-	20	1596847	12+4-	INS	-97	29	2	COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	1600723	3+2-	20	1600747	3+2-	INS	-116	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1608606	6+5-	20	1608612	2+3-	INS	-159	38	5	COLO-829BL-IL|2:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1618061	2+2-	20	1618102	2+2-	INS	-223	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1627702	2+1-	20	1627869	1+2-	INS	-151	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1639749	2+3-	20	1639741	2+3-	INS	-101	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1646680	2+2-	20	1646689	2+2-	INS	-377	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1658457	3+3-	20	1658460	3+3-	INS	-268	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1658825	3+2-	20	1658820	3+2-	INS	-254	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1694600	17+0-	20	1694666	12+30-	DEL	113	99	17	COLO-829BL-IL|4:COLO-829-IL|13	0.44	BreakDancerMax-0.0.1r81	|q10|o20
20	1707810	2+3-	20	1707798	2+3-	INS	-90	32	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1708835	2+2-	20	1708824	2+2-	INS	-238	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1710786	2+2-	20	1710791	2+2-	INS	-238	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1715166	2+2-	20	1715183	2+2-	INS	-103	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1741901	2+3-	20	1741944	2+3-	INS	-248	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1742372	2+0-	20	1742449	0+2-	INS	-244	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1768308	7+1-	20	1768448	1+4-	DEL	138	73	4	COLO-829BL-IL|2:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	1500315	12+1-	20	1850304	14+4-	INV	349909	99	12	COLO-829BL-IL|5:COLO-829-IL|7	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	1768308	3+1-	20	1768784	0+3-	DEL	172	76	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	1770488	4+1-	20	1770563	1+4-	INS	-187	52	5	COLO-829_v2_74|3:COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	1772572	5+4-	20	1772692	5+4-	INS	-292	12	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1775562	2+2-	20	1775574	2+2-	INS	-105	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1781380	2+2-	20	1781367	2+2-	INS	-116	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1782642	2+0-	20	1782781	0+2-	INS	-155	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1796730	12+4-	20	1796832	12+4-	INS	-288	12	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1802759	2+2-	20	1802746	2+2-	INS	-114	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1805768	8+8-	20	1805850	8+8-	INS	-259	54	6	COLO-829_v2_74|4:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	1828591	4+2-	20	1828621	4+2-	INS	-113	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1846449	2+0-	20	1846522	2+3-	INS	-153	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1851970	2+1-	20	1852088	1+2-	INS	-172	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1853323	3+0-	20	1853468	0+2-	INS	-173	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1875176	2+2-	20	1875207	2+2-	INS	-242	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1880298	2+1-	20	1880297	0+2-	INS	-199	25	2	COLO-829_v2_74|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	1896684	3+1-	20	1896753	0+2-	INS	-172	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1897830	2+2-	20	1897835	2+2-	INS	-105	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1900254	4+2-	20	1900281	4+2-	INS	-91	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1901307	2+2-	20	1901338	2+2-	INS	-90	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1923328	5+3-	20	1923360	0+2-	INS	-251	40	5	COLO-829BL-IL|1:COLO-829_v2_74|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	1929615	3+1-	20	1929741	0+2-	INS	-160	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1930281	2+2-	20	1930235	2+2-	INS	-110	40	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1955492	3+1-	20	1955536	0+2-	INS	-268	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	1975951	2+2-	20	1975963	2+2-	INS	-99	29	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	1983873	2+2-	20	1983836	2+2-	INS	-105	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1987038	2+3-	20	1987046	2+3-	INS	-341	19	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	1988389	2+2-	20	1988357	2+2-	INS	-114	36	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2005797	2+0-	20	2005857	3+5-	INS	-211	31	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	2022887	2+2-	20	2022840	2+2-	INS	-397	29	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2029396	2+2-	20	2029344	2+2-	INS	-106	42	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	2060884	2+2-	20	2060824	2+2-	INS	-119	41	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2066629	2+0-	20	2066798	0+4-	INS	-149	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2074264	2+3-	20	2074325	2+3-	INS	-357	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2080481	2+2-	20	2080450	2+2-	INS	-255	26	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2093583	2+2-	20	2093581	2+2-	INS	-93	27	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2094996	5+3-	20	2095007	5+3-	INS	-103	40	3	COLO-829BL-IL|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	2096083	3+2-	20	2096116	3+2-	INS	-252	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2123933	2+2-	20	2123919	2+2-	INS	-117	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	2131549	5+6-	20	2131658	5+6-	INS	-222	39	5	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2140680	2+2-	20	2140714	2+2-	INS	-98	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2142931	5+3-	20	2143013	5+3-	INS	-120	34	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2169707	16+2-	20	2169787	1+15-	DEL	98	99	13	COLO-829BL-IL|4:COLO-829-IL|9	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	2174629	2+2-	20	2174595	2+2-	INS	-115	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2180097	2+0-	20	2180271	0+2-	INS	-150	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2189297	2+0-	20	2189302	0+2-	INS	-194	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2190251	2+2-	20	2190271	2+2-	INS	-213	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2206198	2+2-	20	2206144	2+2-	INS	-116	37	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2210169	3+2-	20	2210161	3+2-	INS	-118	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2222914	2+2-	20	2222940	2+2-	INS	-244	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	2236810	2+0-	20	2236960	0+2-	INS	-178	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2238724	3+5-	20	2238722	3+5-	INS	-274	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2257561	2+2-	20	2257562	2+2-	INS	-246	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	2260664	2+0-	20	2260697	0+3-	INS	-236	16	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2274781	3+0-	20	2274941	1+4-	INS	-238	30	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2292746	3+2-	20	2292782	3+2-	INS	-227	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2295011	2+3-	20	2295050	2+3-	INS	-234	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2307905	15+12-	20	2308601	0+16-	DEL	713	99	13	COLO-829BL-IL|8:COLO-829-IL|5	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	2307905	2+12-	20	2308312	2+0-	ITX	34	55	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2307905	2+10-	20	2308478	12+0-	ITX	509	99	10	COLO-829BL-IL|2:COLO-829-IL|8	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2308610	2+0-	20	2308601	0+3-	INS	-220	12	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	2358018	3+3-	20	2358009	3+3-	INS	-111	45	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2358186	2+2-	20	2358158	2+2-	INS	-108	35	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2395519	2+1-	20	2395597	1+2-	INS	-213	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2400546	2+3-	20	2400619	2+3-	INS	-231	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2413274	3+1-	20	2413299	0+2-	INS	-223	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2436722	2+0-	20	2436736	1+3-	INS	-182	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	2439528	2+2-	20	2439493	2+2-	INS	-90	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2447909	3+0-	20	2448025	0+3-	INS	-205	38	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2471163	3+1-	20	2471223	0+3-	INS	-264	35	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2501535	2+0-	20	2501587	0+2-	INS	-272	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2503723	2+2-	20	2503722	2+2-	INS	-104	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2506925	2+3-	20	2506936	2+3-	INS	-104	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2522827	2+2-	20	2522859	2+2-	INS	-233	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2532688	2+2-	20	2532706	2+2-	INS	-228	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	2535829	2+2-	20	2535813	2+2-	INS	-96	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2540113	2+0-	20	2540101	0+2-	INS	-328	20	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2557409	11+2-	20	2557440	11+2-	INS	-120	24	2	COLO-829-IL|2	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	2565000	2+2-	20	2564992	2+2-	INS	-233	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2578634	2+2-	20	2578672	2+2-	INS	-202	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2583586	2+0-	20	2583630	0+2-	INS	-277	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2592201	3+0-	20	2592252	1+2-	INS	-240	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2618643	2+2-	20	2618620	2+2-	INS	-373	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2628467	3+1-	20	2628558	0+4-	INS	-194	28	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2633814	2+2-	20	2633833	2+2-	INS	-98	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2635511	3+4-	20	2635527	3+4-	INS	-377	30	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2653718	2+2-	20	2653714	2+2-	INS	-239	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2686970	2+2-	20	2686929	2+2-	INS	-109	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2691551	3+0-	20	2691741	0+3-	INS	-135	25	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2693652	2+2-	20	2693662	3+2-	INS	-286	15	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2695444	2+2-	20	2695402	2+2-	INS	-115	34	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	2697421	2+2-	20	2697410	2+2-	INS	-237	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2707308	2+2-	20	2707279	2+2-	INS	-96	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	2744762	2+2-	20	2744755	2+2-	INS	-104	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2751202	39+2-	20	2754408	1+38-	DEL	3265	99	36	COLO-829BL-IL|13:COLO-829-IL|23	0.68	BreakDancerMax-0.0.1r81	|q10|o20
20	2755518	2+0-	20	2755652	0+2-	INS	-186	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2758541	2+2-	20	2758514	2+2-	INS	-94	35	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2771500	11+11-	20	2771539	11+11-	INS	-98	99	11	COLO-829BL-IL|2:COLO-829-IL|9	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	2772612	3+4-	20	2772699	3+4-	INS	-162	24	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2777483	5+3-	20	2777604	5+3-	INS	-99	17	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2807603	2+2-	20	2807588	2+2-	INS	-88	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2809185	2+2-	20	2809205	2+2-	INS	-240	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2812016	25+0-	20	2812325	2+31-	DEL	327	99	24	COLO-829BL-IL|6:COLO-829-IL|18	0.33	BreakDancerMax-0.0.1r81	|q10|o20
20	2844480	5+3-	20	2844528	5+3-	INS	-287	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2847363	3+3-	20	2847380	3+3-	INS	-90	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	2852673	2+0-	20	2852794	0+3-	INS	-181	17	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2867057	2+2-	20	2867027	2+2-	INS	-120	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2874448	2+3-	20	2874412	2+3-	INS	-113	37	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	2875779	2+3-	20	2875813	2+3-	INS	-108	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2883137	2+2-	20	2883119	2+2-	INS	-113	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2898271	17+0-	20	2898366	0+18-	DEL	109	99	17	COLO-829BL-IL|9:COLO-829-IL|8	0.81	BreakDancerMax-0.0.1r81	|q10|o20
20	2911834	2+2-	20	2911783	2+2-	INS	-400	30	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2954339	2+2-	20	2954300	2+2-	INS	-98	37	2	COLO-829BL-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	2963667	2+2-	20	2963635	2+2-	INS	-251	25	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	2969063	3+0-	20	2969269	0+2-	INS	-125	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2969788	22+0-	20	2970076	0+18-	DEL	298	99	17	COLO-829BL-IL|5:COLO-829-IL|12	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	2969788	5+0-	20	2970377	0+3-	DEL	306	73	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	2972723	2+3-	20	2972743	2+3-	INS	-373	17	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	2978537	2+2-	20	2978520	2+2-	INS	-103	29	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	2985948	23+1-	20	2986428	1+2-	DEL	309	43	2	COLO-829_v2_74|2	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	2985948	21+1-	20	2986187	1+21-	DEL	320	99	20	COLO-829BL-IL|7:COLO-829-IL|13	0.56	BreakDancerMax-0.0.1r81	|q10|o20
20	3041374	2+5-	20	3041366	2+5-	INS	-383	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3045269	2+3-	20	3045291	2+3-	INS	-228	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3064779	3+2-	20	3064822	3+2-	INS	-373	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3073223	2+2-	20	3073185	2+2-	INS	-388	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3077038	2+2-	20	3077089	2+2-	INS	-88	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	3078918	3+0-	20	3078942	1+2-	INS	-275	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3079623	2+3-	20	3079643	2+3-	INS	-92	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3087527	2+1-	20	3087617	0+2-	INS	-221	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3103763	2+2-	20	3103761	2+2-	INS	-90	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3128256	3+0-	20	3128336	0+4-	INS	-228	29	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	3205952	2+2-	20	3205993	2+2-	INS	-350	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3218853	2+0-	20	3218930	0+2-	INS	-238	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3248637	2+2-	20	3248629	2+2-	INS	-106	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	3261925	2+2-	20	3261896	2+2-	INS	-86	35	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	3262775	2+2-	20	3262787	2+2-	INS	-109	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3267710	3+0-	20	3267725	0+3-	INS	-292	31	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	3268172	2+1-	20	3268272	1+3-	INS	-185	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3293144	3+5-	20	3293195	3+5-	INS	-185	27	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3295686	3+2-	20	3295696	3+2-	INS	-214	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3295819	2+3-	20	3295833	2+3-	INS	-112	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3310504	2+2-	20	3310528	2+2-	INS	-358	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3313077	2+2-	20	3313116	2+2-	INS	-231	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3314633	2+2-	20	3314637	2+2-	INS	-97	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	3353164	4+3-	20	3353179	4+3-	INS	-108	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3358358	2+2-	20	3358361	2+2-	INS	-104	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	3367052	2+2-	20	3367023	2+2-	INS	-96	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	3373317	2+2-	20	3373293	2+2-	INS	-107	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3406224	2+0-	20	3406320	3+4-	INS	-108	19	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	3408554	3+1-	20	3408661	1+2-	INS	-156	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3430165	3+1-	20	3430217	0+2-	INS	-283	29	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3433631	2+0-	20	3433731	2+2-	INS	-187	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3434916	5+3-	20	3434945	5+3-	INS	-252	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	3437244	3+4-	20	3437269	3+4-	INS	-99	38	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3437679	2+0-	20	3437738	0+2-	INS	-244	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3474292	3+5-	20	3474378	3+5-	INS	-112	30	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3486232	3+3-	20	3486298	3+3-	INS	-107	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	3489399	2+2-	20	3489356	2+2-	INS	-105	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3489749	3+2-	20	3489739	3+2-	INS	-88	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3491854	2+0-	20	3491851	2+4-	INS	-140	39	4	COLO-829_v2_74|1:COLO-829-IL|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	3493030	4+3-	20	3493178	0+2-	INS	-121	27	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3499725	2+3-	20	3499757	2+3-	INS	-382	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3502837	3+2-	20	3502826	3+2-	INS	-109	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3519844	2+0-	20	3519924	1+3-	INS	-204	36	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3532744	2+2-	20	3532768	2+2-	INS	-357	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3541947	3+3-	20	3541977	3+3-	INS	-308	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	3551138	2+0-	20	3551254	0+2-	INS	-215	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3552411	4+5-	20	3552530	4+5-	INS	-257	30	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3568720	2+0-	20	3568872	0+2-	INS	-176	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3570725	2+2-	20	3570682	2+2-	INS	-116	35	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3582117	2+3-	20	3582104	2+3-	INS	-125	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	3595564	2+3-	20	3595628	2+3-	INS	-86	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3596232	4+1-	20	3596391	0+3-	INS	-214	27	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	3596997	2+2-	20	3597012	2+2-	INS	-238	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3625830	3+3-	20	3625890	3+3-	INS	-275	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	3632270	2+2-	20	3632294	2+2-	INS	-96	24	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3687267	2+0-	20	3687281	0+2-	INS	-306	21	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	3692486	2+2-	20	3692440	2+2-	INS	-395	28	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	3695908	2+2-	20	3695918	2+2-	INS	-363	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3745262	3+0-	20	3745332	1+3-	INS	-255	26	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3749624	2+2-	20	3749672	2+2-	INS	-221	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3759270	2+2-	20	3759246	2+2-	INS	-120	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3775084	2+2-	20	3775096	2+2-	INS	-102	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3778320	2+2-	20	3778274	2+2-	INS	-116	36	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3801418	2+4-	20	3801451	2+4-	INS	-98	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3839763	3+2-	20	3839743	3+2-	INS	-87	33	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3856148	2+2-	20	3856135	2+2-	INS	-235	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3858708	2+2-	20	3858678	2+2-	INS	-100	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	3865121	2+2-	20	3865110	2+2-	INS	-101	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3901038	3+2-	20	3901021	3+2-	INS	-400	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3907960	3+2-	20	3907975	3+2-	INS	-106	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	3960510	3+0-	20	3960511	0+4-	INS	-101	50	3	COLO-829BL-IL|1:COLO-829-IL|2	1.00	BreakDancerMax-0.0.1r81	|q10|o20
20	3961065	6+0-	20	3961197	0+4-	DEL	91	95	4	COLO-829BL-IL|2:COLO-829-IL|2	0.67	BreakDancerMax-0.0.1r81	|q10|o20
20	3968963	2+0-	20	3968962	1+4-	INS	-344	20	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	3980466	2+2-	20	3980511	2+2-	INS	-218	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3990774	2+3-	20	3990780	2+3-	INS	-225	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	3993158	2+2-	20	3993151	2+2-	INS	-98	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4020671	3+2-	20	4020748	3+2-	INS	-224	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	4023198	2+2-	20	4023193	2+2-	INS	-102	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4028903	2+1-	20	4029065	0+2-	INS	-160	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4030773	6+29-	20	4030930	6+29-	INS	-94	62	6	COLO-829BL-IL|2:COLO-829-IL|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	4053624	5+5-	20	4053598	5+5-	INS	-87	65	4	COLO-829BL-IL|2:COLO-829-IL|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	4063395	2+0-	20	4063454	0+2-	INS	-270	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4067607	3+9-	20	4067737	3+9-	INS	-100	22	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	4071509	3+2-	20	4071503	3+2-	INS	-355	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4076077	2+2-	20	4076074	2+2-	INS	-108	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4080730	3+0-	20	4080856	0+3-	INS	-164	27	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	4100251	2+2-	20	4100212	2+2-	INS	-389	26	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	4105056	5+2-	20	4105065	0+4-	INS	-252	44	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	4121032	2+2-	20	4121051	2+2-	INS	-220	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4123911	3+3-	20	4123878	3+3-	INS	-308	39	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4150219	2+2-	20	4150226	2+2-	INS	-218	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	4151281	2+2-	20	4151275	2+2-	INS	-94	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	4153167	3+2-	20	4153180	3+2-	INS	-99	25	2	COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	4158549	2+3-	20	4158523	2+3-	INS	-388	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4165096	3+3-	20	4165053	3+3-	INS	-396	44	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4166535	5+7-	20	4166614	5+7-	INS	-365	13	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	4170558	2+0-	20	4170636	0+2-	INS	-247	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4182143	3+0-	20	4182202	0+3-	INS	-257	33	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	4183116	2+2-	20	4183097	2+2-	INS	-99	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	4212098	2+3-	20	4212128	2+3-	INS	-219	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4252000	3+1-	20	4252036	0+2-	INS	-306	34	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	4257411	2+2-	20	4257395	2+2-	INS	-113	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	4292192	4+1-	20	4292239	1+3-	INS	-224	36	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4292514	3+1-	20	4292690	1+2-	INS	-135	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4299770	6+6-	20	4299949	6+6-	INS	-267	33	5	COLO-829_v2_74|4:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4318460	3+3-	20	4318544	3+3-	INS	-108	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4319131	2+2-	20	4319138	2+2-	INS	-102	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	4341128	2+0-	20	4341194	0+2-	INS	-206	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4342048	3+4-	20	4342109	3+4-	INS	-169	26	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4355401	2+2-	20	4355417	2+2-	INS	-106	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4356621	2+4-	20	4356599	2+4-	INS	-110	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4386243	2+2-	20	4386211	2+2-	INS	-115	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4396002	4+3-	20	4396052	4+3-	INS	-178	27	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4396682	3+3-	20	4396709	3+3-	INS	-106	39	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4427913	2+2-	20	4427857	2+2-	INS	-121	40	2	COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	4430421	3+3-	20	4430423	3+3-	INS	-87	30	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4430663	2+1-	20	4430785	1+3-	INS	-150	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4454547	2+0-	20	4454716	2+4-	INS	-133	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4460919	3+3-	20	4460924	3+3-	INS	-295	32	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4470595	2+2-	20	4470599	2+2-	INS	-111	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4486906	2+3-	20	4486936	2+3-	INS	-101	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4534270	2+0-	20	4534303	0+2-	INS	-269	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4538277	3+2-	20	4538278	3+2-	INS	-348	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4544616	2+2-	20	4544584	2+2-	INS	-97	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	4562295	2+2-	20	4562344	2+2-	INS	-236	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4563454	2+0-	20	4563506	0+2-	INS	-286	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4566819	2+3-	20	4566807	2+3-	INS	-93	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4578394	2+2-	20	4578442	2+2-	INS	-194	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	4585499	3+2-	20	4585684	1+2-	INS	-122	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4586662	2+2-	20	4586646	2+2-	INS	-240	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4587258	2+2-	20	4587289	2+2-	INS	-209	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4618946	2+3-	20	4618977	2+3-	INS	-110	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	4620602	2+2-	20	4620573	2+2-	INS	-379	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4624531	2+2-	20	4624510	2+2-	INS	-109	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4629677	2+2-	20	4629659	2+2-	INS	-107	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4630290	2+2-	20	4630256	2+2-	INS	-98	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	4633586	4+2-	20	4633652	4+2-	INS	-105	25	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	4655393	3+2-	20	4655411	3+2-	INS	-373	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4656787	2+3-	20	4656875	2+3-	INS	-89	18	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4657423	2+2-	20	4657388	2+2-	INS	-99	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4662332	2+2-	20	4662313	2+2-	INS	-108	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4664484	3+3-	20	4664514	3+3-	INS	-194	34	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4669955	2+1-	20	4669962	3+3-	INS	-287	13	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4694593	2+4-	20	4694592	2+4-	INS	-123	27	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4699092	2+3-	20	4699175	2+3-	INS	-103	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4704637	2+2-	20	4704675	2+2-	INS	-103	23	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4705362	2+0-	20	4705414	0+3-	INS	-262	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4723395	3+2-	20	4723491	3+2-	INS	-236	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4732375	2+3-	20	4732412	2+3-	INS	-248	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4739852	25+26-	20	4739941	25+26-	INS	-96	99	25	COLO-829BL-IL|5:COLO-829-IL|20	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	4755396	7+0-	20	4756176	1+9-	DEL	755	99	6	COLO-829BL-IL|2:COLO-829-IL|4	0.30	BreakDancerMax-0.0.1r81	|q10|o20
20	4766280	4+4-	20	4766385	4+4-	INS	-369	21	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4783313	2+2-	20	4783305	2+2-	INS	-259	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	4796537	2+2-	20	4796555	2+2-	INS	-94	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4804332	2+1-	20	4804495	1+4-	INS	-127	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	4805543	2+2-	20	4805534	2+2-	INS	-106	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	4808899	2+3-	20	4808952	2+3-	INS	-337	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4822607	4+0-	20	4822603	0+2-	INS	-318	16	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	4832186	2+2-	20	4832162	2+2-	INS	-235	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	4849721	2+3-	20	4849764	2+3-	INS	-99	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4852270	2+0-	20	4852412	0+2-	INS	-173	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4865023	2+0-	20	4865079	0+2-	INS	-267	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4880221	2+2-	20	4880186	2+2-	INS	-107	36	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4887377	3+3-	20	4887405	3+3-	INS	-100	39	3	COLO-829-IL|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	4888974	2+2-	20	4888970	2+2-	INS	-243	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4915715	2+2-	20	4915715	2+2-	INS	-95	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4927707	3+2-	20	4927738	3+2-	INS	-101	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4933094	2+2-	20	4933129	2+2-	INS	-348	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4937721	4+3-	20	4937769	4+3-	INS	-357	26	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4945567	2+2-	20	4945511	2+2-	INS	-406	33	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4961993	2+2-	20	4961970	2+2-	INS	-99	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4971978	3+2-	20	4972036	1+5-	INS	-138	30	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	4981910	2+2-	20	4981884	2+2-	INS	-124	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4988124	2+2-	20	4988091	2+2-	INS	-105	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	4995741	2+3-	20	4995729	2+3-	INS	-396	21	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	5001648	2+3-	20	5001712	2+3-	INS	-96	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5004150	2+1-	20	5004245	0+2-	INS	-231	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5006147	34+1-	20	5006204	1+28-	DEL	132	99	26	COLO-829BL-IL|14:COLO-829-IL|12	0.23	BreakDancerMax-0.0.1r81	|q10|o20
20	5006147	8+1-	20	5006478	0+5-	DEL	128	67	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	5032673	1+1-	20	5032743	2+4-	INS	-110	15	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5033072	2+2-	20	5033023	2+2-	INS	-263	32	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5059851	2+4-	20	5059852	2+4-	INS	-349	19	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5067786	5+2-	20	5067897	1+3-	INS	-229	18	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5079071	4+1-	20	5079116	0+3-	INS	-211	30	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	5080266	5+3-	20	5080287	5+3-	INS	-117	24	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5121196	2+2-	20	5121179	2+2-	INS	-98	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5124014	2+2-	20	5124049	2+2-	INS	-109	23	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5126908	2+2-	20	5126958	2+2-	INS	-106	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5152356	2+3-	20	5152325	2+3-	INS	-102	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5165123	2+2-	20	5165123	2+2-	INS	-99	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5170828	2+2-	20	5170831	2+2-	INS	-248	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5181017	2+2-	20	5181021	2+2-	INS	-364	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5181303	2+2-	20	5181290	2+2-	INS	-252	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5192163	3+2-	20	5192177	3+2-	INS	-112	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5192993	2+2-	20	5192956	2+2-	INS	-112	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5201884	3+0-	20	5201957	0+3-	INS	-242	36	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5203376	2+0-	20	5203534	0+2-	INS	-152	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5208139	2+1-	20	5208318	0+2-	INS	-137	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5208305	2+2-	20	5208264	2+2-	INS	-117	34	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	5210709	2+2-	20	5210711	2+2-	INS	-115	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5223407	3+1-	20	5223444	2+3-	INS	-197	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5235740	2+2-	20	5235715	2+2-	INS	-104	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5257953	3+3-	20	5257974	3+3-	INS	-110	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5260340	3+3-	20	5260336	3+3-	INS	-249	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5261553	2+2-	20	5261528	2+2-	INS	-101	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5261664	2+0-	20	5261762	0+2-	INS	-243	31	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5262038	2+0-	20	5262123	0+2-	INS	-247	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5271325	2+2-	20	5271298	2+2-	INS	-93	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5287304	2+0-	20	5287344	0+2-	INS	-280	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5290456	2+2-	20	5290469	2+2-	INS	-109	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5295868	2+2-	20	5295869	2+2-	INS	-105	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5332594	2+0-	20	5332641	0+2-	INS	-273	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5334245	2+3-	20	5334253	2+3-	INS	-119	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5335700	2+2-	20	5335661	2+2-	INS	-105	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5338215	5+3-	20	5338224	5+3-	INS	-108	39	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5338294	2+0-	20	5338319	1+3-	INS	-272	22	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5358422	2+2-	20	5358441	2+2-	INS	-110	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5363530	2+2-	20	5363496	2+2-	INS	-120	32	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5370009	3+3-	20	5370095	3+3-	INS	-234	15	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5376565	2+2-	20	5376539	2+2-	INS	-119	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5397190	2+0-	20	5397255	0+2-	INS	-263	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5399265	2+2-	20	5399219	2+2-	INS	-396	28	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5406922	2+3-	20	5406894	2+3-	INS	-97	35	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5417301	2+3-	20	5417315	2+3-	INS	-242	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5422764	2+2-	20	5422755	2+2-	INS	-261	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5424359	2+0-	20	5424458	2+5-	INS	-129	22	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5458173	3+0-	20	5458245	2+2-	INS	-250	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5458624	3+2-	20	5458680	6+2-	INS	-220	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5465747	2+2-	20	5465698	2+2-	INS	-113	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	5467461	2+2-	20	5467401	2+2-	INS	-124	41	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5478851	3+0-	20	5478951	0+3-	INS	-237	43	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	5479154	2+2-	20	5479129	2+2-	INS	-99	30	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5530360	3+2-	20	5530405	3+2-	INS	-212	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5531276	2+3-	20	5531264	2+3-	INS	-100	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5550275	2+0-	20	5550360	0+2-	INS	-221	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5570282	2+1-	20	5570268	0+3-	INS	-215	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	5574875	3+1-	20	5575039	0+4-	INS	-167	27	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	5598313	2+2-	20	5598342	2+2-	INS	-221	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5616570	3+1-	20	5616575	1+3-	INS	-294	24	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5620911	4+1-	20	5620903	3+3-	INS	-246	37	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	5622353	3+1-	20	5622384	1+5-	INS	-194	14	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5627887	7+4-	20	5627999	7+4-	INS	-201	12	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5628069	5+2-	20	5628050	5+17-	INS	-121	51	8	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|4	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	5633042	3+2-	20	5632999	3+2-	INS	-114	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5644322	2+2-	20	5644328	2+2-	INS	-109	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5649072	2+2-	20	5649093	2+2-	INS	-238	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5669953	2+0-	20	5670123	2+3-	INS	-151	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5675833	2+3-	20	5675846	2+3-	INS	-103	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5684581	2+2-	20	5684571	2+2-	INS	-239	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5699711	2+2-	20	5699753	2+2-	INS	-102	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5704283	2+0-	20	5704353	0+2-	INS	-259	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5716259	2+3-	20	5716237	2+3-	INS	-241	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5717151	2+0-	20	5717204	0+2-	INS	-277	24	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	5724772	2+1-	20	5724801	0+4-	INS	-235	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5725537	2+2-	20	5725561	2+2-	INS	-100	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5747993	2+2-	20	5748008	2+2-	INS	-241	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5750425	2+2-	20	5750384	2+2-	INS	-111	34	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5767593	2+2-	20	5767582	2+2-	INS	-393	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5769171	2+2-	20	5769160	2+2-	INS	-110	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5776012	2+1-	20	5776080	0+4-	INS	-208	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5780537	3+2-	20	5780518	3+2-	INS	-96	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5808400	2+2-	20	5808429	2+2-	INS	-90	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5834275	2+2-	20	5834234	2+2-	INS	-104	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5843322	3+3-	20	5843372	3+3-	INS	-92	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5871928	2+2-	20	5871947	2+2-	INS	-210	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5875813	2+2-	20	5875859	2+2-	INS	-94	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5908113	2+2-	20	5908148	2+2-	INS	-90	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5912788	2+0-	20	5912905	0+2-	INS	-206	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5915490	2+2-	20	5915474	2+2-	INS	-98	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5926887	4+1-	20	5926958	0+3-	INS	-184	40	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	5943043	3+0-	20	5943200	0+3-	INS	-160	36	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	5975052	2+0-	20	5975134	0+2-	INS	-241	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	5977485	2+1-	20	5977468	2+4-	INS	-260	33	3	COLO-829_v2_74|2:COLO-829-IL|1	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	5983594	2+2-	20	5983550	2+2-	INS	-111	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	5990949	2+1-	20	5990948	2+3-	INS	-241	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	5999858	2+2-	20	5999810	2+2-	INS	-398	29	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6034201	2+0-	20	6034192	1+3-	INS	-253	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	6035207	3+3-	20	6035284	3+3-	INS	-154	24	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6040954	3+1-	20	6041156	0+2-	INS	-112	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6043652	2+2-	20	6043641	2+2-	INS	-109	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	6061106	2+2-	20	6061063	2+2-	INS	-249	29	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6068020	3+1-	20	6068036	1+3-	INS	-282	38	4	COLO-829_v2_74|3:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	6079217	2+2-	20	6079226	2+2-	INS	-91	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6098956	32+0-	20	6099484	0+2-	DEL	325	43	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6098956	30+0-	20	6099276	1+33-	DEL	334	99	30	COLO-829BL-IL|14:COLO-829_v2_74|1:COLO-829-IL|15	0.24	BreakDancerMax-0.0.1r81	|q10|o20
20	6101487	5+3-	20	6101586	5+3-	INS	-178	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6101656	3+1-	20	6101788	0+2-	INS	-159	11	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6106229	2+2-	20	6106302	2+2-	INS	-92	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6108080	2+2-	20	6108089	2+2-	INS	-98	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6118846	2+2-	20	6118813	2+2-	INS	-103	36	2	COLO-829BL-IL|2	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	5310485	0+3-	20	6198314	0+3-	INV	887737	59	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6137936	2+2-	20	6137935	2+2-	INS	-94	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	6169509	2+2-	20	6169508	0+2-	INS	-290	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6187976	2+2-	20	6187980	2+2-	INS	-115	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6199201	5+0-	20	6199294	0+5-	DEL	97	98	5	COLO-829BL-IL|1:COLO-829-IL|4	0.16	BreakDancerMax-0.0.1r81	|q10|o20
20	6220628	3+2-	20	6220722	0+2-	INS	-177	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6222570	3+1-	20	6222651	0+2-	INS	-283	30	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6231346	2+3-	20	6231333	2+3-	INS	-395	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6238324	2+2-	20	6238321	2+2-	INS	-97	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	6255931	2+2-	20	6255881	2+2-	INS	-114	37	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6287332	5+0-	20	6287322	1+6-	INS	-326	65	6	COLO-829_v2_74|6	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	6289619	2+0-	20	6289641	0+2-	INS	-318	30	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6299423	3+0-	20	6299559	0+3-	INS	-181	33	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6310429	3+4-	20	6310418	3+4-	INS	-105	42	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6330647	3+4-	20	6330661	3+4-	INS	-291	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6337702	3+0-	20	6337727	1+3-	INS	-310	41	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	6368991	3+3-	20	6369008	3+3-	INS	-261	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6369937	3+3-	20	6369959	3+3-	INS	-123	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	6378676	2+4-	20	6378828	1+3-	INS	-151	37	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	6381517	2+2-	20	6381482	2+2-	INS	-107	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6401422	2+3-	20	6401412	2+3-	INS	-106	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6420649	2+2-	20	6420638	2+2-	INS	-230	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6424405	2+3-	20	6424377	2+3-	INS	-109	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	6427311	2+2-	20	6427274	2+2-	INS	-93	37	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6429240	2+2-	20	6429238	2+2-	INS	-384	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6435083	2+2-	20	6435068	2+2-	INS	-99	33	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6446688	2+0-	20	6446723	0+2-	INS	-293	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6452319	2+2-	20	6452287	2+2-	INS	-381	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6452808	2+0-	20	6452878	0+2-	INS	-254	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6459062	2+0-	20	6459151	0+2-	INS	-244	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6484867	3+2-	20	6484868	3+2-	INS	-89	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6485065	2+3-	20	6485214	2+3-	INS	-99	17	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6494349	2+0-	20	6494378	0+2-	INS	-273	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6507210	2+2-	20	6507182	2+2-	INS	-378	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6508220	2+2-	20	6508210	2+2-	INS	-103	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6508721	2+3-	20	6508754	2+3-	INS	-94	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	6524425	2+3-	20	6524434	2+3-	INS	-242	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6544883	2+2-	20	6544848	2+2-	INS	-99	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6546443	3+0-	20	6546580	0+2-	INS	-162	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6572492	2+0-	20	6572687	0+2-	INS	-122	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6589353	2+0-	20	6589562	1+3-	INS	-122	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6593814	7+8-	20	6593861	7+8-	INS	-96	98	7	COLO-829BL-IL|1:COLO-829-IL|6	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6608762	2+0-	20	6608883	0+3-	INS	-166	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6620102	2+2-	20	6620077	2+2-	INS	-99	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6638455	2+3-	20	6638450	2+3-	INS	-378	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6638688	2+3-	20	6638692	2+3-	INS	-110	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6646786	2+2-	20	6646796	2+2-	INS	-240	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6653789	2+1-	20	6653864	1+3-	INS	-189	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6668869	2+0-	20	6669050	0+2-	INS	-133	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6670864	3+0-	20	6671042	1+3-	INS	-146	16	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	6687193	2+2-	20	6687173	2+2-	INS	-99	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6695782	2+2-	20	6695803	2+2-	INS	-90	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6697766	2+2-	20	6697787	2+2-	INS	-96	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6704225	2+3-	20	6704311	2+3-	INS	-97	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6712140	2+0-	20	6712220	0+2-	INS	-255	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6743432	4+2-	20	6743414	1+2-	INS	-277	31	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6743777	2+0-	20	6743903	0+2-	INS	-195	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6756575	2+2-	20	6756578	2+2-	INS	-97	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6769915	20+23-	20	6770112	20+23-	INS	-175	99	19	COLO-829BL-IL|1:COLO-829_v2_74|8:COLO-829-IL|10	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	6778836	5+4-	20	6778941	5+4-	INS	-283	12	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6779011	2+2-	20	6779072	0+2-	INS	-172	10	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6793497	6+5-	20	6793632	6+5-	INS	-213	41	5	COLO-829_v2_74|2:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6828581	4+1-	20	6828616	3+3-	INS	-223	26	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	6844651	2+2-	20	6844673	2+2-	INS	-224	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	6851751	10+3-	20	6851898	10+3-	INS	-87	16	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6852725	3+3-	20	6852734	3+3-	INS	-101	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6855415	2+2-	20	6855553	0+2-	INS	-141	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6871242	2+2-	20	6871259	2+2-	INS	-239	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6873232	2+2-	20	6873209	2+2-	INS	-244	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6882423	2+2-	20	6882454	2+2-	INS	-113	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6889223	2+2-	20	6889270	2+2-	INS	-221	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6892329	2+3-	20	6892288	2+3-	INS	-105	38	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6918040	3+2-	20	6918028	3+2-	INS	-361	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6918268	3+4-	20	6918290	3+4-	INS	-110	40	3	COLO-829-IL|3	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	6932494	2+2-	20	6932453	2+2-	INS	-98	38	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6933738	2+0-	20	6933819	0+2-	INS	-241	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6945006	3+2-	20	6945041	0+2-	INS	-224	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6945782	4+4-	20	6945895	4+4-	INS	-207	29	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	6952289	3+3-	20	6952273	3+3-	INS	-241	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	6968772	3+3-	20	6968816	3+3-	INS	-170	27	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	6969716	2+0-	20	6969809	0+2-	INS	-223	16	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	7000547	2+2-	20	7000526	2+2-	INS	-95	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7016043	2+2-	20	7016017	2+2-	INS	-116	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7056096	2+2-	20	7056117	2+2-	INS	-213	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	7073903	2+7-	20	7073965	2+7-	INS	-338	14	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7082374	2+1-	20	7082418	0+2-	INS	-291	24	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	7105490	2+2-	20	7105462	2+2-	INS	-110	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	7106729	2+0-	20	7106794	0+2-	INS	-252	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7118192	3+2-	20	7118259	3+2-	INS	-234	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	7124340	2+3-	20	7124385	2+3-	INS	-219	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7137901	2+2-	20	7137892	2+2-	INS	-105	32	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	7149796	2+2-	20	7149769	2+2-	INS	-110	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7170326	2+0-	20	7170493	0+2-	INS	-151	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7201522	5+4-	20	7201647	5+4-	INS	-283	11	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7204258	3+4-	20	7204276	3+4-	INS	-184	32	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7222085	6+1-	20	7222596	2+66-	DEL	318	99	5	COLO-829_v2_74|5	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	7222347	61+0-	20	7222596	2+61-	DEL	317	99	61	COLO-829BL-IL|19:COLO-829-IL|42	0.73	BreakDancerMax-0.0.1r81	|q10|o20
20	7284607	2+0-	20	7284645	0+2-	INS	-273	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7292708	3+2-	20	7292719	3+2-	INS	-99	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7309100	2+2-	20	7309115	2+2-	INS	-235	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7312562	2+2-	20	7312549	2+2-	INS	-104	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	7315616	2+2-	20	7315611	2+2-	INS	-224	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7322268	3+1-	20	7322356	0+3-	INS	-204	28	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7323726	2+3-	20	7323788	2+3-	INS	-204	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	7329808	2+2-	20	7329775	2+2-	INS	-99	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7393088	3+2-	20	7393152	3+2-	INS	-95	25	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7403784	2+2-	20	7403764	2+2-	INS	-93	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7405783	2+2-	20	7405799	2+2-	INS	-106	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	7408181	2+2-	20	7408145	2+2-	INS	-385	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7423953	3+2-	20	7423952	3+2-	INS	-120	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7444372	2+2-	20	7444348	2+2-	INS	-241	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7454072	2+2-	20	7454056	2+2-	INS	-104	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7459422	2+2-	20	7459391	2+2-	INS	-123	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7494930	2+0-	20	7495131	0+2-	INS	-115	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7508192	2+1-	20	7508327	2+4-	INS	-140	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7517300	2+2-	20	7517257	2+2-	INS	-100	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7537034	2+3-	20	7537016	2+3-	INS	-112	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7627563	2+2-	20	7627536	2+2-	INS	-115	31	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7647687	2+3-	20	7647720	2+3-	INS	-201	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7650768	3+2-	20	7650749	3+2-	INS	-120	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7693996	2+2-	20	7694045	2+2-	INS	-89	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7699743	2+0-	20	7699784	0+2-	INS	-277	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7722664	4+2-	20	7722745	4+2-	INS	-96	20	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7733045	2+3-	20	7733091	2+3-	INS	-224	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	7742694	3+2-	20	7742732	3+2-	INS	-96	27	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7763765	2+2-	20	7763782	2+2-	INS	-114	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7766003	3+3-	20	7766074	3+3-	INS	-96	33	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7770571	3+2-	20	7770651	1+3-	INS	-131	39	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7784990	2+2-	20	7784947	2+2-	INS	-114	39	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	7792841	2+0-	20	7792870	2+2-	INS	-195	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7807985	3+1-	20	7808051	0+2-	INS	-180	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7839795	2+3-	20	7839798	2+3-	INS	-89	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7841004	2+2-	20	7840984	2+2-	INS	-96	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7851728	2+2-	20	7851681	2+2-	INS	-115	36	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7853549	2+2-	20	7853507	2+2-	INS	-104	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7856416	2+0-	20	7856431	1+3-	INS	-223	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	7888775	2+2-	20	7888813	2+2-	INS	-104	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7895012	3+3-	20	7895081	3+3-	INS	-101	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7896359	3+5-	20	7896511	3+5-	INS	-219	17	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7904079	3+2-	20	7904213	2+3-	INS	-115	35	4	COLO-829BL-IL|2:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7912160	2+2-	20	7912190	2+2-	INS	-206	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	7913073	2+0-	20	7913079	0+3-	INS	-255	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7926792	2+2-	20	7926775	2+2-	INS	-87	33	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7934708	3+2-	20	7934685	3+2-	INS	-116	34	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7943084	3+2-	20	7943088	3+2-	INS	-395	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7956386	2+4-	20	7956454	2+4-	INS	-117	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7957301	2+2-	20	7957268	2+2-	INS	-382	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	7959292	4+2-	20	7959399	0+3-	INS	-159	34	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7963315	2+2-	20	7963283	2+2-	INS	-95	32	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	7981703	2+0-	20	7981827	2+3-	INS	-115	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	7991270	3+3-	20	7991291	3+3-	INS	-171	30	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8033561	2+2-	20	8033504	2+2-	INS	-407	33	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8036074	3+2-	20	8036034	3+2-	INS	-107	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8051968	2+3-	20	8052012	2+3-	INS	-105	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8067422	2+2-	20	8067405	2+2-	INS	-108	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8071953	2+2-	20	8071945	2+2-	INS	-231	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8085343	2+3-	20	8085320	2+3-	INS	-108	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8093149	2+2-	20	8093138	2+2-	INS	-101	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8100004	2+0-	20	8100113	0+2-	INS	-177	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8127717	2+0-	20	8127778	0+2-	INS	-271	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8135647	23+0-	20	8135798	1+25-	DEL	194	99	23	COLO-829BL-IL|7:COLO-829-IL|16	0.27	BreakDancerMax-0.0.1r81	|q10|o20
20	8155521	2+2-	20	8155562	2+2-	INS	-89	23	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	8156082	3+3-	20	8156090	3+3-	INS	-106	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8163168	2+3-	20	8163200	2+3-	INS	-101	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8164974	2+2-	20	8165008	2+2-	INS	-92	23	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8169404	2+3-	20	8169457	2+3-	INS	-102	22	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8173919	2+2-	20	8173890	2+2-	INS	-94	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8174393	2+2-	20	8174388	2+2-	INS	-104	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8179986	2+2-	20	8179939	2+2-	INS	-103	40	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8182277	2+3-	20	8182256	2+3-	INS	-117	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8186958	2+2-	20	8186914	2+2-	INS	-394	28	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8197663	2+2-	20	8197650	2+2-	INS	-122	28	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	8199404	2+2-	20	8199374	2+2-	INS	-107	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8200569	2+0-	20	8200631	2+4-	INS	-266	31	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8208408	2+2-	20	8208380	2+2-	INS	-99	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8211771	2+3-	20	8211789	2+3-	INS	-98	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8215732	3+3-	20	8215742	3+3-	INS	-190	32	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8216220	3+0-	20	8216341	0+5-	INS	-221	34	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	8248975	2+3-	20	8248998	2+3-	INS	-106	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8257642	2+0-	20	8257754	0+2-	INS	-210	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8261619	2+2-	20	8261597	2+2-	INS	-244	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8272687	2+6-	20	8272794	2+6-	INS	-239	14	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8292293	3+2-	20	8292420	3+3-	INS	-206	23	4	COLO-829_v2_74|3:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8301502	2+2-	20	8301515	2+2-	INS	-213	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8303734	2+3-	20	8303787	2+3-	INS	-238	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8319235	2+2-	20	8319258	2+2-	INS	-242	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8331942	2+3-	20	8332007	2+3-	INS	-95	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8342017	2+2-	20	8342004	2+2-	INS	-121	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8344386	2+3-	20	8344406	2+3-	INS	-108	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8346498	2+1-	20	8346644	0+2-	INS	-175	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8351059	2+3-	20	8351159	2+3-	INS	-102	19	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8358995	2+1-	20	8359061	1+3-	INS	-220	36	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8399407	2+2-	20	8399411	2+2-	INS	-110	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8400340	2+3-	20	8400346	2+3-	INS	-226	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8403119	2+2-	20	8403086	2+2-	INS	-115	32	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8417942	2+3-	20	8417914	2+3-	INS	-102	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8419051	2+3-	20	8419051	2+3-	INS	-93	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8422344	7+0-	20	8422451	45+33-	ITX	-161	99	22	COLO-829BL-IL|8:COLO-829-IL|14	0.63	BreakDancerMax-0.0.1r81	|q10|o20
20	8422682	20+1-	20	8422708	0+20-	DEL	153	99	19	COLO-829BL-IL|6:COLO-829-IL|13	0.19	BreakDancerMax-0.0.1r81	|q10|o20
20	8425492	3+0-	20	8425644	1+4-	INS	-192	33	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8433069	2+3-	20	8433145	2+3-	INS	-217	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8433861	4+1-	20	8433921	2+5-	INS	-219	49	6	COLO-829BL-IL|1:COLO-829_v2_74|4:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	8441067	2+2-	20	8441062	2+2-	INS	-95	31	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8457120	2+2-	20	8457133	2+2-	INS	-243	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8464475	2+2-	20	8464482	2+2-	INS	-105	30	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8467156	2+2-	20	8467137	2+2-	INS	-237	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8472760	3+1-	20	8472746	1+3-	INS	-207	36	4	COLO-829_v2_74|2:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	8482275	5+3-	20	8482329	5+3-	INS	-283	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8482399	2+0-	20	8482547	0+2-	INS	-159	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8500542	2+2-	20	8500517	2+2-	INS	-251	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8507914	2+2-	20	8507906	2+2-	INS	-115	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8511314	3+3-	20	8511345	3+3-	INS	-256	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8512438	2+5-	20	8512453	2+5-	INS	-124	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8533549	2+2-	20	8533507	2+2-	INS	-391	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8535686	2+2-	20	8535659	2+2-	INS	-108	31	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8542715	4+3-	20	8542763	4+3-	INS	-104	34	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8543694	2+2-	20	8543687	2+2-	INS	-252	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8544259	3+1-	20	8544359	0+2-	INS	-167	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8545045	2+0-	20	8545056	1+2-	INS	-301	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8551977	4+3-	20	8551989	4+3-	INS	-100	41	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8556365	2+4-	20	8556410	2+4-	INS	-236	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8567000	2+0-	20	8567121	0+3-	INS	-163	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8568057	2+4-	20	8568104	2+4-	INS	-92	22	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8608440	2+0-	20	8608547	1+3-	INS	-186	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8615705	3+2-	20	8615716	3+2-	INS	-109	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8625897	2+3-	20	8625904	2+3-	INS	-349	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8636477	2+2-	20	8636527	2+2-	INS	-336	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8644317	2+0-	20	8644472	0+2-	INS	-183	28	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8648646	2+2-	20	8648629	2+2-	INS	-246	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8651178	2+2-	20	8651144	2+2-	INS	-106	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8666393	2+2-	20	8666370	2+2-	INS	-120	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8671210	2+3-	20	8671218	2+3-	INS	-228	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8697830	3+3-	20	8697896	3+3-	INS	-198	27	3	COLO-829_v2_74|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8709184	2+2-	20	8709184	2+2-	INS	-222	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8716054	2+2-	20	8716076	2+2-	INS	-85	28	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8735091	2+2-	20	8735097	2+2-	INS	-101	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8770796	2+2-	20	8770827	2+2-	INS	-94	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8784640	2+2-	20	8784662	2+2-	INS	-102	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8792040	3+1-	20	8792119	2+4-	INS	-179	39	5	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8793027	3+2-	20	8793021	3+2-	INS	-96	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8804775	2+2-	20	8804740	2+2-	INS	-250	27	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8811007	2+2-	20	8811014	2+2-	INS	-99	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8824637	2+2-	20	8824613	2+2-	INS	-106	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8839807	2+2-	20	8839830	2+2-	INS	-101	24	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8852418	3+3-	20	8852451	3+3-	INS	-192	29	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8857169	2+2-	20	8857150	2+2-	INS	-112	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8860461	2+2-	20	8860465	2+2-	INS	-88	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8869327	2+2-	20	8869351	2+2-	INS	-96	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8872696	2+2-	20	8872715	2+2-	INS	-105	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8883188	2+1-	20	8883309	0+2-	INS	-189	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8899184	4+2-	20	8899257	1+3-	INS	-165	47	5	COLO-829_v2_74|2:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8900447	2+3-	20	8900473	2+3-	INS	-102	28	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8910268	2+0-	20	8910368	1+4-	INS	-175	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8918710	3+2-	20	8918662	3+2-	INS	-123	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	8924751	2+3-	20	8924853	2+3-	INS	-168	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8932225	2+2-	20	8932231	2+2-	INS	-111	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8944262	3+0-	20	8944714	0+4-	DEL	156	82	3	COLO-829_v2_74|3	0.33	BreakDancerMax-0.0.1r81	|q10|o20
20	8950504	4+2-	20	8950561	4+2-	INS	-199	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	8965359	3+2-	20	8965383	3+2-	INS	-97	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	8977154	5+4-	20	8978361	1+5-	DEL	1177	91	4	COLO-829BL-IL|2:COLO-829-IL|2	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	8977154	1+4-	20	8978103	5+0-	ITX	779	84	4	COLO-829BL-IL|2:COLO-829-IL|2	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	8977808	2+2-	20	8977757	2+2-	INS	-401	30	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	8988174	2+1-	20	8988311	1+3-	INS	-150	34	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9001555	2+1-	20	9001597	0+2-	INS	-245	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9010554	2+2-	20	9010516	2+2-	INS	-118	33	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9014369	2+0-	20	9014538	2+3-	INS	-139	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9014840	2+2-	20	9014828	2+2-	INS	-108	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9024868	2+2-	20	9024856	2+2-	INS	-100	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9045347	2+3-	20	9045332	2+3-	INS	-102	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9049535	4+4-	20	9049547	4+4-	INS	-290	41	4	COLO-829_v2_74|3:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	9082561	3+1-	20	9082691	0+2-	INS	-246	30	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9084056	4+1-	20	9084103	0+2-	INS	-185	19	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9089371	2+2-	20	9089329	2+2-	INS	-391	27	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9096340	3+3-	20	9096383	3+3-	INS	-89	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9099648	2+2-	20	9099638	2+2-	INS	-241	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9107915	2+2-	20	9107914	2+2-	INS	-234	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9117282	15+8-	20	9117431	0+6-	INS	-130	62	8	COLO-829BL-IL|2:COLO-829_v2_74|4:COLO-829-IL|2	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	9117282	6+3-	20	9117265	4+7-	DEL	104	63	4	COLO-829BL-IL|2:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	9117406	2+1-	20	9117431	0+2-	INS	-270	15	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	9129161	3+2-	20	9129178	3+2-	INS	-94	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9133816	2+2-	20	9133855	2+2-	INS	-348	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9143367	2+0-	20	9143390	0+3-	INS	-288	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9144007	2+2-	20	9144005	2+2-	INS	-362	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9170894	2+2-	20	9170877	2+2-	INS	-235	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9171101	2+0-	20	9171267	1+3-	INS	-124	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9202081	4+1-	20	9202246	1+2-	INS	-135	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9202914	2+3-	20	9202914	2+3-	INS	-115	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9209244	2+2-	20	9209254	2+2-	INS	-246	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9216574	2+2-	20	9216545	2+2-	INS	-102	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9217202	2+2-	20	9217199	2+2-	INS	-107	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9223830	3+3-	20	9223905	3+3-	INS	-90	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9232893	2+2-	20	9232846	2+2-	INS	-113	36	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9262762	3+1-	20	9262818	1+1-	INS	-190	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9273983	2+2-	20	9273969	2+2-	INS	-89	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9283687	2+2-	20	9283632	2+2-	INS	-115	38	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9296037	2+2-	20	9296042	2+2-	INS	-244	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9307893	2+3-	20	9307934	2+3-	INS	-232	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9314057	4+4-	20	9314047	4+4-	INS	-97	42	3	COLO-829BL-IL|1:COLO-829-IL|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	9327532	2+2-	20	9327523	2+2-	INS	-100	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9334801	2+2-	20	9334814	2+2-	INS	-254	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9355063	2+2-	20	9355055	2+2-	INS	-109	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9364040	3+1-	20	9364046	1+3-	INS	-270	41	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	9398230	2+0-	20	9398330	1+2-	INS	-213	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9405030	2+3-	20	9404996	2+3-	INS	-121	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9410119	2+2-	20	9410133	2+2-	INS	-223	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9414529	2+1-	20	9414533	0+2-	INS	-335	23	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	9434011	3+0-	20	9434049	0+3-	INS	-290	38	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	9460313	2+3-	20	9460330	2+3-	INS	-109	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9467292	2+2-	20	9467260	2+2-	INS	-96	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9470758	2+2-	20	9470703	2+2-	INS	-117	38	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9476636	2+2-	20	9476673	2+2-	INS	-204	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9495835	3+0-	20	9495986	0+4-	INS	-178	33	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	9500696	3+0-	20	9500756	0+2-	INS	-269	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9507643	2+2-	20	9507629	2+2-	INS	-111	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9524204	2+0-	20	9524391	0+2-	INS	-138	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9525849	4+4-	20	9525883	4+4-	INS	-297	38	4	COLO-829_v2_74|3:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9560001	2+2-	20	9559978	2+2-	INS	-88	34	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9581000	2+3-	20	9581022	2+3-	INS	-98	28	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9588980	3+1-	20	9588980	0+8-	INS	-286	11	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	9602278	2+2-	20	9602239	2+2-	INS	-113	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9603333	3+4-	20	9603433	3+4-	INS	-216	20	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9606488	2+2-	20	9606512	2+2-	INS	-100	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9609993	3+3-	20	9609993	3+3-	INS	-198	35	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9617093	3+0-	20	9617184	0+2-	INS	-205	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9618411	4+5-	20	9618553	4+5-	INS	-347	29	4	COLO-829_v2_74|4	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9619987	2+2-	20	9619960	2+2-	INS	-377	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9634799	3+0-	20	9634823	0+3-	INS	-268	30	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	9644787	2+0-	20	9644902	0+2-	DEL	85	42	2	COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	9651795	2+0-	20	9651930	2+4-	INS	-240	25	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9668068	2+2-	20	9668023	2+2-	INS	-105	39	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9670705	3+1-	20	9670698	0+2-	INS	-233	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	9671681	4+0-	20	9671665	0+2-	INS	-213	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	9689137	3+4-	20	9689174	3+4-	INS	-182	30	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9696065	2+2-	20	9696034	2+2-	INS	-98	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9703218	3+2-	20	9703186	3+2-	INS	-122	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9714874	2+3-	20	9714959	2+3-	INS	-299	13	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9719570	2+1-	20	9719668	0+2-	INS	-217	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9747061	2+2-	20	9747092	2+2-	INS	-102	24	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9755680	3+3-	20	9755731	3+3-	INS	-101	26	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9763676	2+2-	20	9763627	2+2-	INS	-125	37	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9766157	2+2-	20	9766175	2+2-	INS	-94	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9766469	2+0-	20	9766596	1+3-	INS	-158	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9768028	2+2-	20	9768022	2+2-	INS	-252	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9837360	2+2-	20	9837379	2+2-	INS	-207	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9855237	2+2-	20	9855209	2+2-	INS	-246	26	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9859740	3+2-	20	9859769	3+2-	INS	-96	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9866914	2+0-	20	9866975	0+3-	INS	-237	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9869983	2+3-	20	9869998	2+3-	INS	-113	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9872233	2+2-	20	9872217	2+2-	INS	-114	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9907315	2+3-	20	9907270	2+3-	INS	-395	28	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	9924979	3+3-	20	9924982	3+3-	INS	-106	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9925331	4+1-	20	9925365	0+4-	INS	-254	36	4	COLO-829_v2_74|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	9952491	2+2-	20	9952509	2+2-	INS	-102	29	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9962220	2+4-	20	9962224	2+4-	INS	-97	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9966006	3+4-	20	9966059	3+4-	INS	-162	28	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9968032	2+3-	20	9968010	2+3-	INS	-99	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9969966	2+2-	20	9969970	2+2-	INS	-104	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9981910	3+2-	20	9981919	3+2-	INS	-104	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9983382	2+2-	20	9983418	2+2-	INS	-202	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	9984489	3+3-	20	9984512	3+3-	INS	-380	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	9989459	2+1-	20	9989457	1+3-	INS	-241	30	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	10008255	2+1-	20	10008366	1+4-	INS	-166	20	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	10010169	2+2-	20	10010163	2+2-	INS	-95	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10011429	3+1-	20	10011499	1+3-	INS	-152	31	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	10017546	3+2-	20	10017638	0+2-	INS	-178	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10021704	2+2-	20	10021693	2+2-	INS	-102	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10035322	2+0-	20	10035418	1+3-	INS	-171	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10048154	6+4-	20	10048170	0+2-	INS	-174	49	6	COLO-829_v2_74|3:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10078751	2+0-	20	10078864	0+2-	DEL	86	41	2	COLO-829-IL|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	10084355	2+2-	20	10084304	2+2-	INS	-401	30	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10138337	2+0-	20	10138484	0+2-	INS	-172	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10166009	2+0-	20	10166093	0+2-	INS	-237	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10177867	2+0-	20	10178058	1+2-	INS	-116	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10180933	2+2-	20	10180895	2+2-	INS	-387	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10190735	2+2-	20	10190709	2+2-	INS	-103	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10193028	2+3-	20	10193034	2+3-	INS	-121	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10199504	2+3-	20	10199519	1+2-	INS	-264	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10203575	2+3-	20	10203610	2+3-	INS	-98	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10209909	2+2-	20	10209927	2+2-	INS	-248	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10221361	2+0-	20	10221584	0+2-	INS	-112	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10222108	3+1-	20	10222112	3+5-	INS	-197	34	4	COLO-829_v2_74|2:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	10232432	2+2-	20	10232416	2+2-	INS	-245	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10252402	2+0-	20	10252461	65+62-	ITX	-144	99	30	COLO-829BL-IL|12:COLO-829-IL|18	0.24	BreakDancerMax-0.0.1r81	|q10|o20
20	10252852	9+4-	20	10252843	0+9-	INS	-143	63	9	COLO-829_v2_74|9	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	10254736	2+1-	20	10254798	1+4-	INS	-238	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10256110	3+2-	20	10256140	3+2-	INS	-236	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10258144	2+2-	20	10258179	2+2-	INS	-98	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10261253	2+1-	20	10261249	0+2-	INS	-273	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10279982	2+2-	20	10279949	2+2-	INS	-383	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10297339	2+3-	20	10297319	2+3-	INS	-369	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10312452	2+0-	20	10312604	0+2-	INS	-174	23	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	10327842	3+0-	20	10327986	0+3-	INS	-172	35	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10365410	2+2-	20	10365390	2+2-	INS	-87	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10385963	2+2-	20	10385947	2+2-	INS	-114	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10388825	2+2-	20	10388846	2+2-	INS	-99	24	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10397102	3+1-	20	10397149	1+3-	INS	-204	57	4	COLO-829_v2_74|2:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	10401047	2+2-	20	10401012	2+2-	INS	-110	32	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	10411070	2+2-	20	10411034	2+2-	INS	-110	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10444417	2+2-	20	10444416	2+2-	INS	-231	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10445299	2+2-	20	10445274	2+2-	INS	-244	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10477579	3+2-	20	10477564	3+2-	INS	-100	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10484233	2+0-	20	10484309	0+2-	INS	-258	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10488741	2+2-	20	10488753	2+2-	INS	-220	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10506140	2+2-	20	10506152	2+2-	INS	-91	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10522713	3+1-	20	10522772	0+3-	INS	-211	24	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10532143	2+0-	20	10532238	0+2-	INS	-218	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10552349	2+3-	20	10552386	2+3-	INS	-102	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10552842	3+2-	20	10552849	3+2-	INS	-102	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10555960	2+3-	20	10555939	2+3-	INS	-370	22	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10560118	2+0-	20	10560287	0+2-	INS	-168	28	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10561301	2+2-	20	10561275	2+2-	INS	-254	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10567343	2+2-	20	10567294	2+2-	INS	-258	30	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10569300	3+3-	20	10569337	3+3-	INS	-103	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10574374	3+3-	20	10574475	0+2-	INS	-124	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10585614	2+2-	20	10585650	2+2-	INS	-94	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10612657	2+2-	20	10612677	2+2-	INS	-104	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10613573	4+2-	20	10613707	0+3-	INS	-122	39	4	COLO-829_v2_74|2:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	10617569	2+1-	20	10617757	0+3-	INS	-125	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10619790	3+1-	20	10619926	0+2-	INS	-154	35	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10622442	2+0-	20	10622498	0+2-	INS	-265	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10627976	2+2-	20	10627962	2+2-	INS	-109	33	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10634227	2+4-	20	10634274	2+4-	INS	-209	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10637642	2+2-	20	10637686	2+2-	INS	-89	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10641297	2+3-	20	10641289	2+3-	INS	-103	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10702443	3+1-	20	10702454	1+2-	INS	-218	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	10708966	3+1-	20	10709100	1+3-	INS	-135	39	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10718391	3+0-	20	10718531	0+2-	INS	-170	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10728707	3+1-	20	10728750	1+3-	INS	-313	32	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10730551	2+2-	20	10730572	2+2-	INS	-96	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10746867	2+2-	20	10746836	2+2-	INS	-115	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10747942	2+4-	20	10747921	2+4-	INS	-96	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10753947	2+2-	20	10753956	2+2-	INS	-229	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10757640	3+2-	20	10757658	3+2-	INS	-104	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10762371	2+0-	20	10762479	0+2-	INS	-213	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10778048	2+2-	20	10778019	2+2-	INS	-106	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10778196	2+2-	20	10778153	2+2-	INS	-114	35	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10800780	2+2-	20	10800734	2+2-	INS	-116	36	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10801762	2+2-	20	10801761	2+2-	INS	-122	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10819504	2+2-	20	10819482	2+2-	INS	-372	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10832258	2+2-	20	10832271	2+2-	INS	-223	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10838214	2+1-	20	10838250	0+2-	INS	-254	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10839786	2+2-	20	10839737	2+2-	INS	-120	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	10839878	2+2-	20	10839884	2+2-	INS	-107	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10842863	3+1-	20	10842847	1+3-	INS	-270	36	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	10848158	2+2-	20	10848128	2+2-	INS	-100	35	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10848941	2+0-	20	10848973	0+3-	INS	-268	18	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	10850433	2+3-	20	10850508	2+3-	INS	-88	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10852958	2+2-	20	10852986	2+2-	INS	-234	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10853749	2+2-	20	10853785	2+2-	INS	-106	27	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10857086	2+2-	20	10857083	2+2-	INS	-97	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10884624	3+0-	20	10884748	0+3-	INS	-176	29	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10892047	2+1-	20	10892110	2+4-	INS	-184	23	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	10902966	3+5-	20	10903045	3+5-	INS	-266	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10904593	2+2-	20	10904573	2+2-	INS	-369	22	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10930377	2+2-	20	10930373	2+2-	INS	-98	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10934795	2+2-	20	10934790	2+2-	INS	-97	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10946683	3+1-	20	10946759	0+2-	INS	-140	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10964298	2+2-	20	10964345	2+2-	INS	-195	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10967450	2+3-	20	10967488	2+3-	INS	-96	27	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10971873	3+4-	20	10971957	3+4-	INS	-284	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	10972725	2+2-	20	10972683	2+2-	INS	-123	34	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	10984781	2+2-	20	10984750	2+2-	INS	-93	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11019330	2+2-	20	11019310	2+2-	INS	-107	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11025839	2+2-	20	11025876	2+2-	INS	-93	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11026276	3+4-	20	11026329	3+4-	INS	-293	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11027093	2+2-	20	11027102	2+2-	INS	-106	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11031549	2+0-	20	11031632	0+2-	INS	-224	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11036405	3+3-	20	11036401	3+3-	INS	-242	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11037213	2+1-	20	11037266	0+2-	INS	-209	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11044426	2+2-	20	11044429	2+2-	INS	-360	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11051054	2+2-	20	11051005	2+2-	INS	-112	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	11064897	2+0-	20	11065026	1+2-	INS	-187	16	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	11065592	2+3-	20	11065615	2+3-	INS	-238	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11084204	2+1-	20	11084232	0+3-	INS	-288	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11092798	2+2-	20	11092801	2+2-	INS	-108	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11096968	2+2-	20	11096929	2+2-	INS	-261	28	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11106695	3+3-	20	11106752	3+3-	INS	-97	35	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11106966	2+2-	20	11106934	2+2-	INS	-95	36	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11108712	2+0-	20	11108895	0+2-	INS	-130	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11122121	4+4-	20	11122187	4+4-	INS	-279	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11133301	2+0-	20	11133293	0+2-	INS	-322	21	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	11135225	2+0-	20	11135213	2+4-	INS	-204	41	4	COLO-829BL-IL|2:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	11151167	2+2-	20	11151108	2+2-	INS	-118	40	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11157678	2+2-	20	11157656	2+2-	INS	-113	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11172505	4+2-	20	11172531	0+2-	INS	-255	25	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11181672	2+2-	20	11181643	2+2-	INS	-103	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11187485	3+2-	20	11187491	3+2-	INS	-95	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11207843	3+3-	20	11207862	3+3-	INS	-227	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11232650	3+1-	20	11232718	0+2-	INS	-182	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11243766	2+2-	20	11243734	2+2-	INS	-381	24	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11253142	2+4-	20	11253169	2+4-	INS	-217	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11255298	2+2-	20	11255301	2+2-	INS	-255	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11270277	2+2-	20	11270301	2+2-	INS	-97	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11270494	3+1-	20	11270490	0+2-	INS	-265	33	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	11273200	2+5-	20	11273177	2+5-	INS	-91	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11276261	3+3-	20	11276256	3+3-	INS	-112	43	3	COLO-829BL-IL|2:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11277561	2+2-	20	11277523	2+2-	INS	-98	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11282530	2+3-	20	11282556	2+3-	INS	-94	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11309423	3+2-	20	11309414	3+2-	INS	-369	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11341374	2+2-	20	11341334	2+2-	INS	-105	34	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	11341977	2+0-	20	11342056	0+2-	INS	-253	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11349622	4+2-	20	11349643	4+2-	INS	-219	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11366315	2+2-	20	11366309	2+2-	INS	-115	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11373080	2+2-	20	11373049	2+2-	INS	-96	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11380400	2+2-	20	11380484	2+2-	INS	-328	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11399213	2+3-	20	11399267	2+3-	INS	-106	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11402626	2+2-	20	11402649	2+2-	INS	-100	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11423240	2+3-	20	11423241	2+3-	INS	-245	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11425591	2+2-	20	11425617	2+2-	INS	-108	24	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11431752	2+2-	20	11431740	2+2-	INS	-116	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11452461	2+0-	20	11452669	0+2-	INS	-112	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11455655	2+3-	20	11455729	2+3-	INS	-239	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11462946	0+2-	20	11466869	0+4-	INV	3854	50	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11465276	93+0-	20	11465867	0+3-	DEL	312	59	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11465276	90+0-	20	11465587	0+83-	DEL	323	99	83	COLO-829BL-IL|20:COLO-829_v2_74|11:COLO-829-IL|52	0.23	BreakDancerMax-0.0.1r81	|q10|o20
20	11465276	7+0-	20	11465763	0+6-	DEL	323	99	6	COLO-829_v2_74|6	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11471216	2+4-	20	11471241	2+4-	INS	-119	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11488752	2+2-	20	11488791	2+2-	INS	-250	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11489551	2+3-	20	11489521	2+3-	INS	-101	35	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11508168	2+2-	20	11508163	2+2-	INS	-113	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11543534	4+4-	20	11543516	4+4-	INS	-246	50	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	11548213	2+2-	20	11548194	2+2-	INS	-259	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11550169	3+2-	20	11550157	3+2-	INS	-101	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11574447	2+2-	20	11574429	2+2-	INS	-92	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11588910	2+0-	20	11588924	2+4-	INS	-313	33	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11595139	2+0-	20	11596676	0+29-	DEL	1245	47	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	11595447	31+0-	20	11596676	0+27-	DEL	1246	99	26	COLO-829BL-IL|9:COLO-829-IL|17	0.17	BreakDancerMax-0.0.1r81	|q10|o20
20	11595447	5+0-	20	11596882	0+5-	DEL	1243	99	5	COLO-829_v2_74|5	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	11631305	2+3-	20	11631325	2+3-	INS	-89	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11631887	3+1-	20	11631990	2+3-	INS	-160	24	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11635133	2+2-	20	11635094	2+2-	INS	-112	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11639919	2+0-	20	11640034	0+2-	INS	-205	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11645966	2+3-	20	11646012	2+3-	INS	-241	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11667109	2+2-	20	11667104	2+2-	INS	-230	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11677691	2+0-	20	11677722	2+3-	INS	-158	20	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11683243	2+0-	20	11683293	0+2-	INS	-258	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11699116	2+9-	20	11699154	2+9-	INS	-352	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11714181	2+1-	20	11714308	0+3-	INS	-214	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11716581	2+0-	20	11716586	0+2-	INS	-309	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11719491	2+4-	20	11719446	2+4-	INS	-108	39	2	COLO-829BL-IL|2	0.33	BreakDancerMax-0.0.1r81	|q10|o20
20	11721362	3+4-	20	11721462	3+4-	INS	-196	24	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11727570	2+2-	20	11727603	2+2-	INS	-93	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11765559	2+3-	20	11765528	2+3-	INS	-96	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11801177	2+3-	20	11801175	2+3-	INS	-231	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11807729	2+2-	20	11807711	2+2-	INS	-108	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11838283	3+2-	20	11838342	1+3-	INS	-222	32	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11874011	2+2-	20	11873972	2+2-	INS	-389	26	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	11886658	3+3-	20	11886702	3+3-	INS	-107	34	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	11904046	3+3-	20	11904093	3+3-	INS	-107	34	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11915557	2+2-	20	11915543	2+2-	INS	-228	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11927535	2+1-	20	11927746	0+2-	INS	-130	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11928637	2+2-	20	11928613	2+2-	INS	-104	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11936913	2+2-	20	11936892	2+2-	INS	-370	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11956939	3+4-	20	11957042	3+4-	INS	-214	14	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11960543	2+3-	20	11960547	2+3-	INS	-124	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11979276	3+2-	20	11979279	3+2-	INS	-98	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11987449	2+2-	20	11987491	2+2-	INS	-91	23	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	11991685	2+2-	20	11991659	2+2-	INS	-110	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11996157	2+2-	20	11996207	2+2-	INS	-233	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	11998863	3+0-	20	11998874	1+3-	INS	-303	14	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	12029305	2+2-	20	12029297	0+2-	INS	-357	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12031953	2+2-	20	12031926	2+2-	INS	-253	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12037649	4+2-	20	12037676	4+2-	INS	-373	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12044459	3+2-	20	12044502	3+2-	INS	-90	27	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12064641	2+2-	20	12064679	2+2-	INS	-97	23	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	12071352	2+2-	20	12071317	2+2-	INS	-98	36	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	12098266	2+2-	20	12098214	2+2-	INS	-117	36	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12111050	3+3-	20	12111083	0+3-	INS	-190	27	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	12113012	2+3-	20	12113027	2+3-	INS	-102	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12126608	2+0-	20	12126648	0+2-	INS	-284	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12129319	4+0-	20	12129452	1+3-	INS	-172	24	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12134745	2+2-	20	12134740	2+2-	INS	-115	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12152554	2+2-	20	12152538	2+2-	INS	-230	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12173607	4+4-	20	12173685	4+4-	INS	-163	38	4	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12181066	2+2-	20	12181085	2+2-	INS	-89	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12189560	2+2-	20	12189526	2+2-	INS	-109	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12194884	3+0-	20	12195012	0+3-	INS	-197	37	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	12213735	2+1-	20	12213818	0+3-	INS	-216	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12216896	3+3-	20	12216941	3+3-	INS	-108	34	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12228821	2+2-	20	12228839	2+2-	INS	-92	29	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12229310	2+3-	20	12229293	2+3-	INS	-92	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12236178	2+3-	20	12236180	2+3-	INS	-98	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12238527	2+2-	20	12238512	2+2-	INS	-100	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	12242286	2+2-	20	12242251	2+2-	INS	-95	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12279500	2+2-	20	12279459	2+2-	INS	-103	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12280092	2+2-	20	12280091	2+2-	INS	-232	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12281687	2+1-	20	12281720	1+3-	INS	-216	32	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12313853	3+3-	20	12313880	3+3-	INS	-105	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12335779	2+2-	20	12335793	2+2-	INS	-210	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	12343883	2+0-	20	12344033	0+2-	INS	-171	21	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	12363715	2+2-	20	12363661	2+2-	INS	-126	39	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	12366413	2+2-	20	12366374	2+2-	ITX	-123	53	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12368610	3+1-	20	12368592	1+2-	INS	-267	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	12368959	2+2-	20	12368977	2+2-	INS	-107	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	12396553	2+1-	20	12396744	0+2-	INS	-115	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12401700	11+12-	20	12401779	11+12-	INS	-90	99	11	COLO-829BL-IL|6:COLO-829-IL|5	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12354468	0+7-	20	12423390	0+7-	INV	68829	99	5	COLO-829-IL|5	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	12427772	2+2-	20	12427730	2+2-	INS	-252	29	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12430846	2+2-	20	12430890	2+2-	INS	-242	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12444595	2+0-	20	12444583	0+2-	INS	-205	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	12450110	3+3-	20	12450158	3+3-	INS	-185	28	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12460898	3+1-	20	12460883	2+5-	INS	-293	47	5	COLO-829_v2_74|5	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	12475327	2+2-	20	12475301	2+2-	INS	-89	35	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12476459	2+0-	20	12476636	0+2-	INS	-144	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12482133	2+2-	20	12482126	2+2-	INS	-87	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12487462	11+9-	20	12487540	11+9-	INS	-96	75	6	COLO-829BL-IL|1:COLO-829-IL|5	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12493408	4+4-	20	12493463	4+4-	INS	-222	41	4	COLO-829BL-IL|2:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12501059	2+1-	20	12501095	0+2-	INS	-298	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12504710	3+4-	20	12504758	3+4-	INS	-188	27	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12538205	2+1-	20	12538222	1+3-	INS	-200	24	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12542051	2+2-	20	12542042	2+2-	INS	-236	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	12562388	3+2-	20	12562407	3+2-	INS	-106	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12574924	2+0-	20	12575104	1+3-	INS	-233	33	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12578583	2+2-	20	12578607	2+2-	INS	-208	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12598554	2+0-	20	12598666	0+2-	INS	-191	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12600754	2+1-	20	12600926	0+2-	INS	-135	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12610813	2+3-	20	12610787	2+3-	INS	-99	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12614590	2+2-	20	12614566	2+2-	INS	-240	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	12620530	2+1-	20	12620549	0+2-	INS	-296	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12623119	2+2-	20	12623083	2+2-	ITX	-129	46	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12626368	2+2-	20	12626349	2+2-	INS	-112	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	12634804	3+3-	20	12634801	3+3-	INS	-197	35	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12637041	2+0-	20	12637231	1+2-	INS	-138	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12657918	2+3-	20	12657938	2+3-	INS	-104	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12663125	4+5-	20	12663200	4+5-	INS	-250	38	4	COLO-829BL-IL|2:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12671994	2+2-	20	12672070	1+3-	INS	-146	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12675932	2+3-	20	12675909	2+3-	INS	-98	34	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12689843	2+2-	20	12689855	2+2-	INS	-94	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	12701911	3+2-	20	12701974	3+2-	INS	-198	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12705067	2+2-	20	12705052	2+2-	INS	-120	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12723585	2+2-	20	12723553	2+2-	INS	-108	36	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12725076	3+2-	20	12725037	3+2-	INS	-403	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12739430	3+2-	20	12739414	3+2-	INS	-112	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	12743270	2+1-	20	12743363	0+2-	INS	-191	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12765940	2+2-	20	12765894	2+2-	ITX	-126	49	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12770530	3+3-	20	12770560	3+3-	INS	-245	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12773121	2+0-	20	12773204	1+3-	INS	-162	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12815690	2+3-	20	12815670	2+3-	INS	-373	22	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	12823818	2+0-	20	12823810	0+2-	INS	-316	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12846757	3+2-	20	12846748	3+2-	INS	-88	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12878264	2+0-	20	12878267	0+2-	INS	-301	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12881606	3+2-	20	12881593	3+2-	INS	-115	28	2	COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	12887927	2+0-	20	12887936	0+3-	INS	-317	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12896883	3+0-	20	12896875	1+3-	INS	-219	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	12905122	3+2-	20	12905181	0+2-	INS	-196	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12908353	3+3-	20	12908363	3+3-	INS	-281	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12914072	2+1-	20	12914115	2+5-	INS	-168	29	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12927599	11+6-	20	12927642	11+6-	ITX	-185	99	6	COLO-829BL-IL|3:COLO-829-IL|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	12927712	5+0-	20	12927811	0+5-	DEL	193	70	4	COLO-829BL-IL|2:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	12930866	3+3-	20	12930896	3+3-	INS	-291	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	12935465	2+2-	20	12935471	2+2-	INS	-96	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12958087	2+2-	20	12958064	2+2-	INS	-104	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12958703	2+2-	20	12958708	2+2-	INS	-94	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12966069	2+0-	20	12966125	0+3-	INS	-248	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	12973957	2+2-	20	12973986	2+2-	INS	-94	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13008832	2+2-	20	13008837	2+2-	INS	-245	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13015787	3+1-	20	13015884	0+4-	INS	-234	33	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13027423	2+3-	20	13027455	2+3-	INS	-98	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13054572	4+1-	20	13054560	0+2-	INS	-244	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13063620	3+1-	20	13063675	1+2-	INS	-192	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13071042	2+3-	20	13071087	2+3-	INS	-91	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13076266	2+2-	20	13076221	2+2-	INS	-119	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13100871	2+2-	20	13100853	2+2-	INS	-96	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13108735	23+1-	20	13112095	0+24-	DEL	3381	99	21	COLO-829-IL|21	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	13108735	2+1-	20	13112333	1+2-	DEL	3357	44	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13130967	2+2-	20	13130912	2+2-	INS	-125	39	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13131441	3+1-	20	13131509	0+2-	INS	-208	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13137120	3+0-	20	13137192	0+3-	INS	-270	39	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13137674	2+2-	20	13137663	2+2-	INS	-97	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13140886	2+3-	20	13140852	2+3-	INS	-383	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13143783	2+1-	20	13143913	0+2-	INS	-172	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13158165	3+1-	20	13158179	0+2-	INS	-164	20	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13173484	2+2-	20	13173456	2+2-	INS	-94	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13174055	2+3-	20	13174136	2+3-	INS	-178	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13179024	2+2-	20	13178998	2+2-	INS	-103	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13183800	2+2-	20	13183797	2+2-	INS	-112	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13188643	2+3-	20	13188624	2+3-	INS	-94	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13190936	3+2-	20	13190936	3+2-	INS	-388	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13192661	2+2-	20	13192654	2+2-	INS	-107	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13193717	2+3-	20	13193691	2+3-	INS	-105	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13212522	2+2-	20	13212495	2+2-	INS	-112	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13214821	2+2-	20	13214827	2+2-	INS	-105	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13225181	3+0-	20	13225295	0+3-	INS	-202	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13234786	2+0-	20	13234911	0+2-	INS	-199	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13269557	2+2-	20	13269530	2+2-	INS	-376	23	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13273070	2+0-	20	13273160	0+2-	INS	-234	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13281558	2+3-	20	13281592	2+3-	INS	-221	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13284671	2+2-	20	13284660	2+2-	INS	-384	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13298182	2+2-	20	13298162	2+2-	INS	-109	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13312392	2+2-	20	13312399	2+2-	INS	-94	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13322106	2+2-	20	13322127	2+2-	INS	-249	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13337861	2+3-	20	13337837	2+3-	INS	-112	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13340035	2+0-	20	13340082	1+3-	INS	-265	20	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	13354700	2+2-	20	13354650	2+2-	INS	-125	37	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13370257	2+4-	20	13370253	2+4-	ITX	-131	41	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13378907	3+3-	20	13378944	3+3-	INS	-188	33	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13405843	2+2-	20	13405819	2+2-	INS	-251	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13434802	2+2-	20	13434766	2+2-	INS	-386	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13436074	3+2-	20	13436116	3+2-	INS	-97	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13470163	2+0-	20	13470239	0+2-	INS	-261	28	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13497250	2+2-	20	13497220	2+2-	INS	-98	35	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13499092	2+1-	20	13499204	0+2-	INS	-181	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13516166	2+4-	20	13516258	2+4-	INS	-194	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13517160	2+1-	20	13517253	0+2-	INS	-220	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13534975	2+2-	20	13534923	2+2-	INS	-115	36	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13561583	2+3-	20	13561567	2+3-	INS	-110	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13567037	2+3-	20	13567068	2+3-	INS	-348	16	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13571141	2+0-	20	13571276	0+2-	INS	-195	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13587511	2+2-	20	13587560	2+2-	INS	-100	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13600670	3+2-	20	13600661	3+2-	INS	-241	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13612248	2+0-	20	13612365	0+2-	INS	-195	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13620372	2+1-	20	13620450	0+2-	INS	-247	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13621098	2+0-	20	13621222	1+4-	INS	-130	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13627106	2+2-	20	13627081	2+2-	INS	-375	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13665945	2+2-	20	13665915	2+2-	INS	-253	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13695525	3+4-	20	13695531	3+4-	INS	-99	39	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13708529	2+3-	20	13708552	2+3-	INS	-102	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13711014	2+2-	20	13710997	2+2-	INS	-106	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	13716313	2+2-	20	13716295	2+2-	INS	-368	22	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	13716926	2+2-	20	13716918	2+2-	INS	-119	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13728469	2+3-	20	13728484	2+3-	INS	-97	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13733490	2+2-	20	13733470	2+2-	INS	-94	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13733979	4+6-	20	13734069	4+6-	INS	-101	47	4	COLO-829-IL|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13748658	2+2-	20	13748630	2+2-	INS	-378	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13753987	2+2-	20	13753994	2+2-	INS	-376	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13755245	2+2-	20	13755257	2+2-	INS	-217	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13761290	2+2-	20	13761294	2+2-	INS	-104	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13775921	2+2-	20	13775883	2+2-	INS	-102	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13777172	12+2-	20	13777153	8+4-	ITX	-129	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	13777172	10+0-	20	13777345	2+4-	INS	-222	24	4	COLO-829_v2_74|4	0.20	BreakDancerMax-0.0.1r81	|q10|o20
20	13777888	2+2-	20	13777867	2+2-	INS	-401	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13790613	2+2-	20	13790587	2+2-	INS	-242	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13793414	2+3-	20	13793452	2+3-	INS	-106	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13803347	2+0-	20	13803411	0+2-	INS	-257	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13834371	6+3-	20	13834402	6+3-	INS	-93	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13842380	2+2-	20	13842333	2+2-	ITX	-131	50	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13863113	16+5-	20	13863095	0+10-	INS	-98	99	9	COLO-829BL-IL|4:COLO-829-IL|5	0.60	BreakDancerMax-0.0.1r81	|q10|o20
20	13864295	4+4-	20	13864403	4+4-	INS	-142	35	4	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13865642	3+1-	20	13865626	2+3-	INS	-147	38	4	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	13868607	2+2-	20	13868595	0+3-	INS	-91	30	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	13868914	3+2-	20	13868887	3+2-	INS	-111	35	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13920137	2+1-	20	13920155	0+3-	INS	-319	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13935905	2+3-	20	13935867	2+3-	INS	-269	26	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13967042	2+4-	20	13967076	2+4-	INS	-108	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13968771	2+2-	20	13968760	2+2-	INS	-111	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13977680	2+2-	20	13977703	2+2-	INS	-245	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	13982676	3+3-	20	13982732	3+3-	INS	-98	35	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	13994610	2+3-	20	13994616	2+3-	INS	-109	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	14000728	3+1-	20	14000894	8+3-	INS	-132	21	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14001068	8+1-	20	14001138	1+10-	DEL	94	99	8	COLO-829BL-IL|1:COLO-829-IL|7	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	14004009	3+1-	20	14004023	0+2-	INS	-221	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14013058	2+3-	20	14013032	2+3-	INS	-253	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	14046825	2+2-	20	14046804	2+2-	INS	-106	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14048168	2+1-	20	14048218	0+3-	INS	-278	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14079707	2+0-	20	14079709	1+3-	INS	-300	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14081551	4+1-	20	14081596	0+4-	INS	-217	38	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	14086917	2+2-	20	14086862	2+2-	INS	-117	39	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	14091792	3+2-	20	14091828	3+2-	INS	-229	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14103712	2+3-	20	14103701	2+3-	INS	-237	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14111636	4+0-	20	14111662	4+3-	INV	-78	99	4	COLO-829BL-IL|1:COLO-829-IL|3	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	14111751	0+3-	20	14111821	0+3-	INV	-41	94	3	COLO-829-IL|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	14112924	2+2-	20	14112897	2+2-	INS	-112	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14113310	3+3-	20	14113368	3+3-	INS	-224	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14116584	2+2-	20	14116533	2+2-	INS	-122	38	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14127076	3+4-	20	14127183	3+4-	INS	-108	29	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14133126	2+0-	20	14133233	0+2-	INS	-226	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14133805	2+2-	20	14133806	2+2-	INS	-246	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14145092	5+2-	20	14145110	5+2-	INS	-95	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14148187	3+2-	20	14148243	3+2-	INS	-100	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14149792	3+0-	20	14149797	1+4-	INS	-171	40	4	COLO-829_v2_74|2:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	14162460	2+6-	20	14162491	2+6-	INS	-98	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	14166069	2+2-	20	14166084	2+2-	INS	-240	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	14168598	2+3-	20	14168591	2+3-	INS	-93	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14173039	2+2-	20	14173050	2+2-	INS	-220	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14173602	2+4-	20	14173611	2+4-	INS	-92	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14188824	2+2-	20	14188816	2+2-	INS	-110	32	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14208193	2+3-	20	14208305	2+3-	INS	-218	12	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14222262	2+3-	20	14222264	2+3-	INS	-116	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14224639	2+2-	20	14224597	2+2-	INS	-99	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14227277	3+3-	20	14227299	3+3-	INS	-101	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	14242666	2+2-	20	14242666	2+2-	INS	-229	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14247644	2+0-	20	14247693	0+2-	INS	-281	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14248717	2+2-	20	14248687	2+2-	INS	-100	35	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14251386	3+0-	20	14251393	1+2-	INS	-308	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14256965	2+2-	20	14256946	2+2-	INS	-125	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14259323	2+2-	20	14259328	2+2-	INS	-102	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14262742	2+3-	20	14262802	2+3-	INS	-93	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14267872	5+2-	20	14267896	0+3-	INS	-210	32	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14268149	2+2-	20	14268116	2+2-	INS	-100	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14273518	3+2-	20	14273534	3+2-	INS	-96	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14285777	2+2-	20	14285748	2+2-	INS	-242	26	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	14293498	2+2-	20	14293468	2+2-	INS	-95	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14294881	2+0-	20	14294894	1+2-	INS	-301	21	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	14300681	2+2-	20	14300677	2+2-	INS	-99	31	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	14346398	2+3-	20	14346411	2+3-	INS	-121	29	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14360418	2+3-	20	14360426	2+3-	INS	-103	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14374857	2+2-	20	14374845	2+2-	INS	-238	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14377004	2+3-	20	14377019	2+3-	INS	-95	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14381658	2+0-	20	14381828	0+2-	INS	-148	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14416802	2+2-	20	14416770	2+2-	INS	-93	36	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14420279	2+0-	20	14420389	0+2-	INS	-190	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14439346	2+0-	20	14439468	0+2-	INS	-194	20	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	14440937	2+2-	20	14440911	2+2-	INS	-404	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14448442	2+4-	20	14448488	2+4-	INS	-101	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14477137	59+2-	20	14477638	0+7-	DEL	315	99	7	COLO-829_v2_74|7	0.17	BreakDancerMax-0.0.1r81	|q10|o20
20	14477137	51+1-	20	14477374	0+47-	DEL	316	99	47	COLO-829BL-IL|8:COLO-829-IL|39	0.57	BreakDancerMax-0.0.1r81	|q10|o20
20	14477137	4+1-	20	14477773	0+3-	DEL	332	69	3	COLO-829_v2_74|3	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	14479287	3+1-	20	14479355	1+3-	INS	-264	34	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	14489031	3+3-	20	14489022	3+3-	INS	-290	33	3	COLO-829_v2_74|2:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	14506443	2+0-	20	14506641	0+2-	INS	-133	25	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	14512685	2+2-	20	14512676	2+2-	INS	-111	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14519795	12+18-	20	14521846	3+12-	DEL	2069	99	12	COLO-829BL-IL|2:COLO-829-IL|10	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14519795	0+18-	20	14521556	19+1-	ITX	1677	99	18	COLO-829BL-IL|5:COLO-829-IL|13	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	14522081	3+0-	20	14522125	0+3-	INS	-230	18	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14556440	2+2-	20	14556446	2+2-	INS	-109	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14557118	2+1-	20	14557272	1+2-	INS	-151	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14558394	2+2-	20	14558390	2+2-	INS	-109	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14579086	3+4-	20	14579203	3+4-	INS	-244	19	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14581895	2+2-	20	14581866	2+2-	INS	-91	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	14582847	2+2-	20	14582786	2+2-	ITX	-128	57	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14595672	2+2-	20	14595675	2+2-	INS	-101	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14596560	2+2-	20	14596524	2+2-	INS	-107	33	2	COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	14601955	3+3-	20	14601950	3+3-	INS	-124	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14602776	2+5-	20	14602776	3+5-	INS	-196	27	4	COLO-829_v2_74|2:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	14614322	2+2-	20	14614287	2+2-	INS	-109	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14629153	4+3-	20	14629122	4+3-	INS	-398	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14639561	2+2-	20	14639521	2+2-	INS	-389	26	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	14676254	2+2-	20	14676269	2+2-	INS	-106	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14679904	2+0-	20	14680032	0+2-	INS	-190	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14689650	2+4-	20	14689674	2+4-	INS	-101	24	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	14704788	2+0-	20	14704982	0+2-	INS	-135	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14733485	2+2-	20	14733480	2+2-	INS	-104	31	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	14747382	4+4-	20	14747379	4+4-	INS	-105	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14750539	3+2-	20	14750689	0+2-	INS	-137	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14755484	2+4-	20	14755507	2+4-	INS	-243	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14781526	2+0-	20	14781651	0+2-	INS	-185	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14787100	2+2-	20	14787098	2+2-	INS	-102	31	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	14797440	2+0-	20	14797445	0+2-	INS	-187	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14798447	2+2-	20	14798406	2+2-	INS	-102	38	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14813374	2+2-	20	14813351	2+2-	INS	-107	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14827521	2+2-	20	14827515	2+2-	INS	-114	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	14851467	3+3-	20	14851486	3+3-	INS	-249	30	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14859931	2+0-	20	14860025	0+2-	INS	-228	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14888856	2+0-	20	14888861	0+2-	INS	-189	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	14893769	2+2-	20	14893722	2+2-	INS	-104	40	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14897582	2+2-	20	14897598	2+2-	INS	-95	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14920728	2+2-	20	14920752	2+2-	INS	-247	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14938531	2+2-	20	14938486	2+2-	INS	-118	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14943036	2+0-	20	14943064	1+2-	INS	-288	20	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	14910771	3+0-	20	14962083	0+3-	DEL	51001	51	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	14910996	12+0-	20	14961836	1+18-	DEL	51000	99	9	COLO-829-IL|9	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	14910996	3+0-	20	14962279	0+2-	DEL	50988	47	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14948619	9+0-	20	14961836	1+9-	DEL	13222	99	9	COLO-829-IL|9	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14967337	3+1-	20	14967513	0+2-	INS	-225	29	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	14976404	1+1-	20	14976418	1+4-	INS	-191	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14997029	3+2-	20	14997077	0+2-	INS	-236	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15050636	2+0-	20	15050673	0+2-	INS	-295	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	14936807	3+0-	20	15056818	1+5-	DEL	120003	61	3	COLO-829-IL|3	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	15052456	2+2-	20	15052463	2+2-	INS	-103	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15062062	2+2-	20	15062067	2+2-	INS	-113	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15069882	20+9-	20	15069919	20+9-	INS	-112	98	7	COLO-829BL-IL|3:COLO-829-IL|4	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	15069989	13+2-	20	15070111	0+13-	DEL	103	99	13	COLO-829BL-IL|7:COLO-829-IL|6	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	15075043	3+1-	20	15075063	0+2-	INS	-228	38	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	15093342	2+2-	20	15093307	2+2-	INS	-102	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15093934	3+2-	20	15093949	3+2-	INS	-111	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15118299	2+0-	20	15118351	0+2-	INS	-269	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15148755	2+2-	20	15148761	2+2-	INS	-107	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15157388	3+2-	20	15157425	3+2-	INS	-110	23	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15176569	3+3-	20	15176513	3+3-	INS	-117	60	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15213576	2+2-	20	15213599	2+2-	INS	-94	28	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15222334	2+0-	20	15222373	1+3-	INS	-263	16	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	15249537	5+1-	20	15251765	0+33-	DEL	2030	45	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15249537	3+1-	20	15251925	0+3-	DEL	2058	77	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15249744	30+0-	20	15251765	0+31-	DEL	2034	99	30	COLO-829BL-IL|8:COLO-829_v2_74|1:COLO-829-IL|21	0.23	BreakDancerMax-0.0.1r81	|q10|o20
20	15257059	2+2-	20	15257082	2+2-	INS	-99	24	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15258866	2+2-	20	15258879	2+2-	INS	-110	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15259414	2+2-	20	15259374	2+2-	INS	-266	27	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	15274091	2+2-	20	15274077	2+2-	INS	-101	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15274862	2+2-	20	15274842	2+2-	INS	-245	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15285584	2+2-	20	15285563	2+2-	INS	-370	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15286342	3+3-	20	15286302	3+3-	INS	-103	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	15294978	2+2-	20	15294985	2+2-	INS	-100	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15297539	2+2-	20	15297497	2+2-	INS	-107	34	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15311575	2+2-	20	15311629	2+2-	INS	-236	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15313879	2+3-	20	15313850	2+3-	INS	-250	26	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15330399	2+3-	20	15330397	2+3-	INS	-250	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15344792	2+0-	20	15344947	1+2-	INS	-163	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15346499	2+2-	20	15346508	2+2-	INS	-222	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15375804	2+2-	20	15375768	2+2-	INS	-110	33	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15376219	3+1-	20	15376262	0+2-	INS	-216	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15389251	2+2-	20	15389203	2+2-	INS	-119	36	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15394595	2+1-	20	15394584	1+3-	INS	-93	35	3	COLO-829BL-IL|1:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	15406322	2+2-	20	15406330	2+2-	INS	-108	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15408800	2+2-	20	15408784	2+2-	INS	-112	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15415648	2+2-	20	15415664	2+2-	INS	-93	29	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15417094	4+1-	20	15417234	0+3-	INS	-224	40	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15441750	2+2-	20	15441719	2+2-	INS	-95	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15451461	4+1-	20	15451666	0+2-	INS	-113	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15461644	2+0-	20	15461829	0+2-	INS	-139	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15463425	2+2-	20	15463399	2+2-	INS	-382	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15473924	2+2-	20	15473889	2+2-	INS	-91	36	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15489586	3+3-	20	15489623	3+3-	INS	-94	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15491122	4+4-	20	15491213	4+4-	INS	-174	38	4	COLO-829_v2_74|1:COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15497776	2+2-	20	15497786	2+2-	INS	-107	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15507296	3+3-	20	15507268	3+3-	INS	-91	56	3	COLO-829BL-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15533403	3+1-	20	15533426	1+2-	INS	-227	35	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	15537007	3+1-	20	15537003	1+3-	INS	-234	30	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	15537702	3+1-	20	15537707	1+3-	INS	-262	44	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	15541778	2+2-	20	15541747	2+2-	INS	-381	24	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15547535	2+2-	20	15547491	2+2-	INS	-109	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15550221	2+2-	20	15550194	2+2-	INS	-105	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15551210	2+0-	20	15551373	1+3-	INS	-169	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15562525	2+2-	20	15562526	2+2-	INS	-235	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15582707	2+2-	20	15582672	2+2-	INS	-251	25	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15593425	2+2-	20	15593402	2+2-	INS	-234	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15617344	2+2-	20	15617303	2+2-	INS	-107	38	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15619729	2+2-	20	15619694	2+2-	INS	-109	32	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15632904	2+2-	20	15632912	2+2-	INS	-101	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15633794	2+2-	20	15633749	2+2-	INS	-114	35	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15648856	2+0-	20	15649009	0+3-	INS	-156	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15655142	2+2-	20	15655103	2+2-	INS	-109	33	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15660833	2+3-	20	15660870	2+3-	INS	-108	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15665687	2+2-	20	15665650	2+2-	INS	-104	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15671594	3+2-	20	15671638	0+2-	INS	-250	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15674586	2+2-	20	15674613	2+2-	INS	-245	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15676121	2+2-	20	15676108	2+2-	INS	-107	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15679508	2+1-	20	15679668	0+2-	INS	-110	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15684853	2+2-	20	15684859	2+2-	INS	-104	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15687666	2+2-	20	15687670	2+2-	INS	-94	30	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15695727	2+2-	20	15695748	2+2-	INS	-248	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15699347	3+3-	20	15699337	3+3-	INS	-192	35	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15704814	3+2-	20	15704903	0+2-	INS	-166	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15710082	2+0-	20	15710089	1+2-	INS	-284	17	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	15733919	2+2-	20	15733886	2+2-	INS	-100	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15751916	2+2-	20	15751892	2+2-	INS	-257	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	15774146	2+3-	20	15774162	2+3-	INS	-96	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15790049	3+2-	20	15790038	3+2-	INS	-112	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15796964	3+3-	20	15797031	3+3-	INS	-193	25	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15806838	2+3-	20	15806857	2+3-	INS	-243	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15835437	2+2-	20	15835424	2+2-	INS	-101	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15841585	2+2-	20	15841604	2+2-	INS	-234	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15848409	2+2-	20	15848434	2+2-	INS	-237	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15848703	2+2-	20	15848732	2+2-	INS	-223	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15858614	2+1-	20	15858681	0+2-	INS	-281	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15864628	2+0-	20	15864635	0+2-	INS	-310	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15871035	2+2-	20	15871035	2+2-	INS	-102	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15894533	2+3-	20	15894511	2+3-	INS	-390	23	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15901346	2+2-	20	15901314	2+2-	INS	-110	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15918083	3+3-	20	15918111	3+3-	INS	-108	39	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15925568	2+1-	20	15925727	0+2-	INS	-161	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	15928395	2+2-	20	15928361	2+2-	INS	-99	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15937483	2+2-	20	15937487	2+2-	INS	-105	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15971453	2+2-	20	15971419	2+2-	INS	-96	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	15983603	2+2-	20	15983589	2+2-	INS	-110	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	15994423	2+4-	20	15994431	2+4-	INS	-96	30	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16005336	2+0-	20	16005444	0+3-	INS	-202	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16011350	2+0-	20	16011350	1+3-	INS	-315	25	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	16014701	3+3-	20	16014799	3+3-	INS	-376	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16029914	4+0-	20	16029994	0+5-	INS	-251	41	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16036337	2+3-	20	16036343	2+3-	INS	-104	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16051311	2+2-	20	16051323	2+2-	INS	-107	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16051861	3+0-	20	16051874	1+8-	INS	-207	19	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	16073040	2+2-	20	16072981	2+2-	INS	-127	42	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16082902	2+2-	20	16082868	2+2-	INS	-110	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16089209	2+2-	20	16089242	2+2-	INS	-91	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16106055	2+2-	20	16106049	2+2-	INS	-115	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16117529	118+77-	20	16117511	0+41-	ITX	-14	99	70	COLO-829BL-IL|21:COLO-829_v2_74|13:COLO-829-IL|36	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	16128040	2+0-	20	16128057	0+2-	INS	-188	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	16131418	2+3-	20	16131419	2+3-	INS	-118	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16133996	2+1-	20	16133984	1+4-	INS	-277	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	16144933	2+2-	20	16145066	0+3-	INS	-143	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16148414	2+3-	20	16148422	2+3-	INS	-109	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16158561	2+2-	20	16158544	2+2-	INS	-108	33	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	16162275	3+2-	20	16162299	3+2-	INS	-98	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16168086	2+2-	20	16168030	2+2-	INS	-112	38	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16177525	2+2-	20	16177501	2+2-	INS	-374	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16178379	2+0-	20	16178406	0+2-	INS	-294	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16183107	2+0-	20	16183126	1+3-	INS	-293	27	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	16186587	4+10-	20	16186855	27+4-	ITX	125	99	10	COLO-829BL-IL|2:COLO-829-IL|8	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	16186863	2+7-	20	16186855	19+3-	ITX	-105	99	6	COLO-829BL-IL|3:COLO-829-IL|3	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	16186656	2+2-	20	16186621	2+2-	INS	-107	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16187072	13+1-	20	16187077	0+13-	DEL	90	99	13	COLO-829BL-IL|7:COLO-829-IL|6	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	16201054	2+2-	20	16201062	2+2-	INS	-105	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16204187	2+3-	20	16204175	2+3-	INS	-106	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	16212682	2+0-	20	16212714	0+2-	INS	-267	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16217144	6+8-	20	16217389	3+3-	ITX	-151	57	3	COLO-829BL-IL|1:COLO-829-IL|2	0.21	BreakDancerMax-0.0.1r81	|q10|o20
20	16217144	0+4-	20	16217216	8+2-	ITX	-76	74	4	COLO-829BL-IL|1:COLO-829-IL|3	0.27	BreakDancerMax-0.0.1r81	|q10|o20
20	16217507	3+1-	20	16217505	0+3-	INS	-220	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	16228093	2+2-	20	16228061	2+2-	INS	-99	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16228366	2+0-	20	16228448	0+2-	INS	-229	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16242734	2+0-	20	16242852	1+2-	INS	-192	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16244253	3+3-	20	16244260	3+3-	INS	-300	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16291568	2+3-	20	16291578	2+3-	INS	-95	30	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	16302639	2+2-	20	16302631	2+2-	INS	-100	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16323853	6+2-	20	16324003	0+7-	DEL	142	99	6	COLO-829BL-IL|1:COLO-829-IL|5	0.46	BreakDancerMax-0.0.1r81	|q10|o20
20	16332561	2+3-	20	16332625	2+3-	INS	-101	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16334193	2+2-	20	16334189	2+2-	INS	-93	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16338602	3+0-	20	16338723	2+5-	DEL	100	64	3	COLO-829-IL|3	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	16353306	2+0-	20	16353411	0+2-	INS	-200	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16367192	2+1-	20	16367176	0+2-	INS	-336	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16378543	2+0-	20	16378623	1+4-	INS	-175	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	16387279	2+2-	20	16387254	2+2-	INS	-374	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16444477	2+2-	20	16444428	2+2-	INS	-111	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16455021	2+2-	20	16455029	2+2-	INS	-103	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	16471024	2+2-	20	16471011	2+2-	INS	-95	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16474719	2+1-	20	16474848	0+2-	INS	-188	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16475954	4+2-	20	16476078	0+2-	INS	-141	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16488225	2+0-	20	16488300	1+2-	INS	-261	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16493864	2+0-	20	16493860	4+5-	INS	-192	32	5	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|1	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	16510007	3+1-	20	16509996	1+3-	INS	-240	27	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	16514679	2+2-	20	16514650	2+2-	INS	-259	26	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16517543	3+2-	20	16517603	3+2-	INS	-245	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16538312	3+4-	20	16538393	3+4-	INS	-149	29	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16539790	2+0-	20	16539925	1+3-	INS	-155	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	16544005	2+0-	20	16544108	0+2-	INS	-221	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16553969	3+3-	20	16554066	3+3-	INS	-100	32	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16579918	2+2-	20	16579920	2+2-	INS	-87	30	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16581238	4+3-	20	16581247	4+3-	INS	-201	37	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16589377	3+1-	20	16589464	1+4-	INS	-189	43	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	16595127	2+0-	20	16595267	1+4-	INS	-145	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	16603270	2+2-	20	16603279	2+2-	INS	-233	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16612687	2+2-	20	16612684	2+2-	INS	-108	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	16614963	3+4-	20	16615042	3+4-	INS	-313	23	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16618465	2+0-	20	16618517	1+2-	INS	-257	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16635369	2+3-	20	16635402	2+3-	INS	-115	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16654003	6+3-	20	16654057	6+3-	INS	-295	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16661382	2+0-	20	16661458	1+3-	INS	-199	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16661645	2+2-	20	16661616	2+2-	INS	-106	31	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16664084	3+0-	20	16664211	1+4-	INS	-186	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16665339	2+2-	20	16665304	2+2-	INS	-114	36	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16717728	3+3-	20	16717733	3+3-	INS	-197	32	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16757712	3+3-	20	16757785	3+3-	INS	-99	33	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16758212	2+2-	20	16758179	2+2-	INS	-102	36	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16761351	2+0-	20	16761436	0+2-	INS	-238	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16765274	2+3-	20	16765272	2+3-	INS	-106	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16779570	2+3-	20	16779594	2+3-	INS	-100	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16798790	2+2-	20	16798767	2+2-	INS	-102	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16804111	2+2-	20	16804122	2+2-	INS	-101	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16808486	2+1-	20	16808531	1+3-	INS	-292	24	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16818975	2+2-	20	16818921	2+2-	INS	-403	32	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16836905	2+2-	20	16836847	2+2-	INS	-115	40	2	COLO-829BL-IL|1:COLO-829-IL|1	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	16842961	2+3-	20	16842966	2+3-	INS	-248	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	16845736	2+2-	20	16845714	2+2-	INS	-244	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16856668	2+2-	20	16856625	2+2-	INS	-98	39	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16869209	2+2-	20	16869209	2+2-	INS	-116	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	16872361	4+3-	20	16872446	4+3-	INS	-100	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16875532	4+2-	20	16875596	1+3-	INS	-142	44	5	COLO-829_v2_74|2:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16877240	2+2-	20	16877215	2+2-	INS	-112	34	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16880912	2+3-	20	16880955	2+3-	INS	-91	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16927245	2+0-	20	16927290	0+2-	INS	-277	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16930427	2+2-	20	16930448	2+2-	INS	-219	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16939771	3+1-	20	16939820	0+2-	INS	-223	34	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	16954826	2+3-	20	16954862	2+3-	INS	-95	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	16982160	2+2-	20	16982110	2+2-	INS	-112	37	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	16991150	2+2-	20	16991151	2+2-	INS	-112	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	16991797	2+2-	20	16991748	2+2-	INS	-116	37	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17005755	2+0-	20	17005929	0+3-	INS	-147	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17009948	27+1-	20	17009940	2+24-	DEL	99	99	23	COLO-829BL-IL|2:COLO-829-IL|21	0.35	BreakDancerMax-0.0.1r81	|q10|o20
20	17009948	4+1-	20	17010315	0+4-	DEL	94	92	4	COLO-829_v2_74|4	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	17030553	2+4-	20	17030575	2+4-	INS	-383	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17033717	3+2-	20	17033718	3+2-	INS	-237	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17034244	2+2-	20	17034298	2+2-	INS	-90	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17036849	2+2-	20	17036866	2+2-	INS	-228	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17051237	2+0-	20	17051796	0+38-	DEL	342	45	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	17051511	36+5-	20	17051796	0+36-	DEL	355	99	35	COLO-829BL-IL|14:COLO-829-IL|21	0.92	BreakDancerMax-0.0.1r81	|q10|o20
20	17056100	3+3-	20	17056124	3+3-	INS	-104	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17059931	2+2-	20	17059971	2+2-	INS	-204	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17067227	3+2-	20	17067226	3+2-	INS	-261	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17078381	5+1-	20	17078385	0+3-	INS	-258	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	17078381	2+0-	20	17078579	0+2-	INS	-139	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17086169	2+2-	20	17086127	2+2-	INS	-109	34	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17090210	2+2-	20	17090208	2+2-	INS	-227	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17091205	2+0-	20	17091221	1+2-	INS	-312	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17115733	2+4-	20	17115711	2+4-	INS	-234	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17119385	2+2-	20	17119423	2+2-	INS	-199	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17127498	2+2-	20	17127507	2+2-	INS	-217	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17128688	2+0-	20	17128859	0+2-	INS	-151	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17147664	3+4-	20	17147817	3+4-	INS	-180	11	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17151780	2+3-	20	17151749	2+3-	INS	-101	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17161711	3+3-	20	17161722	3+3-	INS	-112	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17161895	3+0-	20	17161929	0+3-	INS	-296	43	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	17166030	2+3-	20	17166063	2+3-	INS	-212	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17186995	2+3-	20	17187031	2+3-	INS	-100	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17202147	2+0-	20	17202209	0+3-	INS	-243	20	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	17251493	3+2-	20	17251479	3+2-	INS	-92	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17254957	2+3-	20	17254918	2+3-	INS	-107	33	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17261527	2+2-	20	17261535	2+2-	INS	-229	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17264971	2+2-	20	17264920	2+2-	INS	-400	30	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17268789	10+3-	20	17268897	10+3-	INS	-89	31	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17269038	2+7-	20	17269097	2+7-	INS	-111	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17270542	2+1-	20	17270619	0+2-	INS	-216	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17283897	2+2-	20	17283901	2+2-	INS	-106	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17289393	2+2-	20	17289341	2+2-	INS	-122	38	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17305838	2+3-	20	17305869	2+3-	INS	-353	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17313857	2+2-	20	17313972	0+3-	INS	-172	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17321481	2+2-	20	17321516	2+2-	INS	-218	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17327332	2+2-	20	17327448	0+2-	INS	-204	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17328058	2+2-	20	17328062	2+2-	INS	-235	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17328872	2+0-	20	17328878	2+3-	INS	-189	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	17332243	2+2-	20	17332258	2+2-	INS	-104	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17363123	2+2-	20	17363129	2+2-	INS	-91	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17371936	3+3-	20	17371910	3+3-	INS	-288	39	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17378215	2+4-	20	17378228	2+4-	INS	-104	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17388420	2+2-	20	17388391	2+2-	INS	-111	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17389617	2+2-	20	17389628	2+2-	INS	-100	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17392514	2+2-	20	17392496	2+2-	INS	-104	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17393515	3+0-	20	17393517	1+2-	INS	-347	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17400459	2+2-	20	17400477	2+2-	INS	-238	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17445089	2+1-	20	17445163	2+2-	INS	-241	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17445242	2+0-	20	17445234	0+2-	INS	-332	27	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	17448161	2+2-	20	17448162	2+2-	INS	-248	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17454895	2+2-	20	17454902	2+2-	INS	-113	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17467254	2+2-	20	17467241	2+2-	INS	-101	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17470777	3+0-	20	17470953	0+2-	INS	-153	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17479099	2+2-	20	17479043	2+2-	INS	-116	44	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17483330	2+2-	20	17483318	2+2-	INS	-106	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17507713	2+5-	20	17507716	2+5-	INS	-114	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17554889	2+2-	20	17554878	2+2-	INS	-245	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17574278	2+2-	20	17574221	2+2-	INS	-406	33	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17584664	2+0-	20	17584828	0+2-	INS	-155	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17600988	2+2-	20	17600993	2+2-	INS	-94	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17634548	3+0-	20	17634655	0+3-	INS	-226	42	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	17635172	2+2-	20	17635146	2+2-	INS	-110	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17644377	2+2-	20	17644402	2+2-	INS	-245	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17694228	2+2-	20	17694227	0+2-	INS	-349	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17700571	3+1-	20	17700585	0+3-	INS	-273	32	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	17729871	2+2-	20	17729826	2+2-	INS	-110	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17730788	2+3-	20	17730763	2+3-	INS	-94	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17731106	2+0-	20	17731238	0+2-	INS	-187	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17735737	2+2-	20	17735696	2+2-	INS	-106	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17760995	2+2-	20	17760970	2+2-	INS	-249	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17774066	22+1-	20	17774157	0+21-	DEL	115	99	20	COLO-829BL-IL|7:COLO-829-IL|13	0.22	BreakDancerMax-0.0.1r81	|q10|o20
20	17774837	2+3-	20	17774826	2+3-	INS	-265	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17787232	2+1-	20	17787271	2+4-	INS	-252	26	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	17789058	3+1-	20	17789148	1+2-	INS	-201	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17808646	3+0-	20	17808765	0+4-	INS	-199	29	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	17815158	2+2-	20	17815169	2+2-	INS	-109	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	17853848	2+3-	20	17853808	2+3-	INS	-123	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17859168	3+2-	20	17859195	3+2-	INS	-102	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17863151	2+2-	20	17863133	2+2-	INS	-116	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17924115	2+2-	20	17924120	2+2-	INS	-103	26	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	17928193	3+2-	20	17928190	3+2-	INS	-94	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17938008	2+2-	20	17938000	2+2-	INS	-237	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17946872	2+2-	20	17946838	2+2-	INS	-102	36	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17947311	3+3-	20	17947330	3+3-	INS	-276	30	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17950708	7+0-	20	17951354	5+12-	DEL	568	99	7	COLO-829BL-IL|3:COLO-829_v2_74|2:COLO-829-IL|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	17951306	1+4-	20	17951354	5+5-	ITX	-113	88	4	COLO-829-IL|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	17951064	5+0-	20	17951354	1+5-	DEL	307	99	5	COLO-829BL-IL|2:COLO-829-IL|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	17953179	2+2-	20	17953163	2+2-	INS	-96	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	17981529	4+4-	20	17981682	4+4-	INS	-325	19	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17990764	2+2-	20	17990745	2+2-	INS	-98	33	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	17992720	2+2-	20	17992742	2+2-	INS	-90	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18030424	3+3-	20	18030427	3+3-	INS	-97	40	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18040577	2+1-	20	18040863	0+2-	DEL	262	41	2	COLO-829-IL|2	0.50	BreakDancerMax-0.0.1r81	|q10|o20
20	18051425	3+0-	20	18051512	1+2-	INS	-232	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18085227	3+1-	20	18085350	1+3-	INS	-146	21	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18088064	2+2-	20	18088050	2+2-	INS	-110	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18097119	2+2-	20	18097094	2+2-	INS	-119	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18097522	3+3-	20	18097549	3+3-	INS	-105	36	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18100539	3+2-	20	18100542	3+2-	INS	-107	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18109546	2+5-	20	18109582	2+5-	INS	-97	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18135795	2+0-	20	18135895	0+2-	INS	-217	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18138285	86+59-	20	18138336	44+48-	DEL	199	99	53	COLO-829BL-IL|13:COLO-829_v2_74|4:COLO-829-IL|36	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	18138285	8+4-	20	18139244	0+21-	DEL	901	99	6	COLO-829_v2_74|6	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18138285	2+4-	20	18138983	6+2-	ITX	791	63	4	COLO-829BL-IL|4	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18138698	19+0-	20	18138773	0+2-	DEL	89	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18138698	17+0-	20	18139244	0+15-	DEL	576	99	15	COLO-829BL-IL|8:COLO-829-IL|7	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	18138698	2+0-	20	18138890	0+4-	DEL	436	32	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18138989	0+2-	20	18138983	2+0-	ITX	-161	40	2	COLO-829BL-IL|1:COLO-829-IL|1	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	18148066	2+2-	20	18148052	2+2-	INS	-105	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18179052	2+2-	20	18179051	2+2-	INS	-108	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18184192	2+2-	20	18184196	2+2-	INS	-98	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18198565	2+3-	20	18198612	2+3-	INS	-208	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18203387	3+3-	20	18203415	3+3-	INS	-98	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18222490	4+3-	20	18222491	4+3-	INS	-201	39	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18226311	2+3-	20	18226325	2+3-	INS	-373	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18238609	2+2-	20	18238609	2+2-	INS	-216	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18252814	2+2-	20	18252777	2+2-	INS	-116	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18259840	2+2-	20	18259828	2+2-	INS	-229	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18260953	3+2-	20	18261016	3+2-	INS	-213	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	17708082	3+0-	20	18304002	4+4-	INV	595846	75	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18269864	2+2-	20	18269899	2+2-	INS	-207	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18290028	2+2-	20	18290018	2+2-	INS	-89	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18318967	3+1-	20	18318990	0+2-	INS	-316	30	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18331636	2+3-	20	18331709	2+3-	INS	-188	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18341320	2+1-	20	18341381	1+2-	INS	-266	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18361742	2+3-	20	18361747	2+3-	INS	-98	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18381967	3+3-	20	18381992	3+3-	INS	-191	31	3	COLO-829_v2_74|1:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	18390900	2+2-	20	18390887	2+2-	INS	-93	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18405976	2+2-	20	18405990	2+2-	INS	-93	29	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18426059	2+2-	20	18426126	2+2-	INS	-111	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18428875	3+3-	20	18428856	3+3-	INS	-191	37	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18430624	4+2-	20	18430652	4+2-	INS	-101	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18430722	2+0-	20	18430763	0+2-	INS	-233	12	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18431782	3+3-	20	18431770	3+3-	INS	-297	35	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	18435335	2+0-	20	18435388	0+2-	INS	-273	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18440153	2+2-	20	18440139	2+2-	INS	-99	33	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18455985	2+2-	20	18456020	2+2-	INS	-88	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18456919	2+3-	20	18456910	2+3-	INS	-106	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18460622	2+0-	20	18460682	0+3-	INS	-274	27	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	18483555	2+2-	20	18483578	2+2-	INS	-235	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18513076	3+2-	20	18513160	3+2-	INS	-353	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18266901	2+0-	20	18534739	3+2-	DEL	267823	43	2	COLO-829BL-IL|1:COLO-829-IL|1	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	18524242	2+2-	20	18524242	2+2-	INS	-101	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18526492	3+1-	20	18526495	1+2-	INS	-240	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	18540003	0+2-	20	18543821	1+2-	INV	3447	75	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18541932	2+3-	20	18541942	2+3-	INS	-339	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18562930	2+2-	20	18562934	2+2-	INS	-223	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18582803	3+2-	20	18582797	3+2-	INS	-233	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18593041	2+2-	20	18593049	2+2-	INS	-101	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18604583	21+19-	20	18604612	0+2-	INS	-123	99	20	COLO-829BL-IL|7:COLO-829_v2_74|3:COLO-829-IL|10	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	18609618	2+1-	20	18609714	0+2-	INS	-213	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18612820	4+4-	20	18612940	4+4-	INS	-88	17	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18617275	2+2-	20	18617302	2+2-	INS	-98	28	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18618567	23+1-	20	18618631	1+26-	DEL	90	99	23	COLO-829BL-IL|7:COLO-829-IL|16	0.16	BreakDancerMax-0.0.1r81	|q10|o20
20	18624123	12+14-	20	18624169	12+14-	INS	-99	99	12	COLO-829BL-IL|5:COLO-829-IL|7	0.27	BreakDancerMax-0.0.1r81	|q10|o20
20	18679509	2+2-	20	18679489	2+2-	INS	-370	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18681279	2+2-	20	18681286	2+2-	INS	-225	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18696167	2+0-	20	18696172	0+2-	INS	-197	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18696954	3+2-	20	18696977	3+2-	INS	-240	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18708126	2+2-	20	18708150	2+2-	INS	-211	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18712271	2+1-	20	18712384	0+2-	INS	-216	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18732211	2+1-	20	18732268	1+3-	INS	-190	30	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	18749551	2+3-	20	18749553	2+3-	INS	-95	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18754981	3+2-	20	18754963	3+2-	INS	-374	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18756320	2+3-	20	18756404	2+3-	INS	-198	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18776834	2+1-	20	18776900	0+2-	INS	-282	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18778142	3+4-	20	18778169	3+4-	INS	-231	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18813909	3+1-	20	18813967	2+4-	INS	-238	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18815987	3+2-	20	18816053	3+2-	INS	-205	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18824887	2+0-	20	18824998	1+3-	INS	-184	38	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18828496	2+3-	20	18828520	2+3-	INS	-387	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18835726	3+0-	20	18835746	1+2-	INS	-298	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18843499	2+2-	20	18843471	2+2-	INS	-105	35	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18846308	2+1-	20	18846393	0+2-	INS	-196	14	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18851266	2+1-	20	18851373	1+4-	INS	-158	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18851977	3+2-	20	18851939	3+2-	INS	-98	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18852118	2+2-	20	18852153	2+2-	INS	-97	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18853778	3+3-	20	18853775	3+3-	INS	-106	43	3	COLO-829BL-IL|2:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18855987	2+1-	20	18856100	0+2-	INS	-205	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18875847	2+1-	20	18875839	0+2-	INS	-230	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18889508	2+2-	20	18889499	2+2-	INS	-99	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18910682	2+0-	20	18910692	0+2-	INS	-308	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18915174	2+3-	20	18915148	2+3-	INS	-105	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18924824	3+2-	20	18924859	3+2-	INS	-103	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18933345	2+0-	20	18933554	0+2-	INS	-120	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	18952479	3+2-	20	18952551	3+2-	INS	-189	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	18957152	3+3-	20	18957187	3+3-	INS	-110	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	18974136	2+3-	20	18974113	2+3-	INS	-114	30	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18978291	2+2-	20	18978285	2+2-	INS	-110	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	18982348	3+1-	20	18982445	0+2-	INS	-285	29	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19009431	41+1-	20	19009725	3+39-	DEL	322	99	39	COLO-829BL-IL|14:COLO-829-IL|25	0.36	BreakDancerMax-0.0.1r81	|q10|o20
20	19009431	2+1-	20	19009933	0+5-	DEL	317	43	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	19009892	3+0-	20	19009933	0+3-	INS	-224	24	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19011702	2+0-	20	19011749	1+4-	INS	-281	26	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	19033101	2+2-	20	19033091	2+2-	INS	-110	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19035147	2+2-	20	19035179	0+2-	INS	-265	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19035533	2+2-	20	19035516	2+2-	INS	-108	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19040324	3+0-	20	19040394	0+3-	INS	-211	25	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19046246	3+3-	20	19046264	3+3-	INS	-98	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19048990	2+3-	20	19049049	2+3-	INS	-196	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19054378	2+0-	20	19054499	3+7-	INS	-108	45	4	COLO-829_v2_74|1:COLO-829-IL|3	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	19060067	2+2-	20	19060082	2+2-	INS	-103	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19067328	2+0-	20	19067403	0+2-	INS	-264	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19074745	2+2-	20	19074716	2+2-	INS	-99	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19079958	2+2-	20	19079952	2+2-	INS	-99	27	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19083503	26+0-	20	19083913	0+3-	DEL	78	46	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	19083503	24+0-	20	19083593	0+15-	DEL	90	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	19127750	2+1-	20	19127764	1+3-	INS	-300	23	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	19134495	2+2-	20	19134513	2+2-	INS	-226	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19144114	2+2-	20	19144088	2+2-	INS	-103	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19197756	2+2-	20	19197810	2+2-	INS	-87	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19201622	3+2-	20	19201602	3+2-	INS	-97	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19213823	2+3-	20	19213811	2+3-	INS	-362	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19222424	2+3-	20	19222454	2+3-	INS	-98	24	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19235949	2+0-	20	19236011	1+3-	INS	-179	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	19245408	2+2-	20	19245413	2+2-	INS	-98	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19257378	2+0-	20	19257481	0+2-	INS	-212	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19262516	2+3-	20	19262594	2+3-	INS	-108	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19274988	4+2-	20	19275069	0+3-	DEL	110	55	3	COLO-829BL-IL|1:COLO-829-IL|2	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	19294611	2+2-	20	19294604	2+2-	INS	-106	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19300663	2+3-	20	19300701	2+3-	INS	-230	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19321961	2+3-	20	19321959	2+3-	INS	-90	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19333446	3+2-	20	19333464	3+2-	INS	-241	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19333780	2+2-	20	19333791	2+2-	INS	-108	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19334944	2+2-	20	19334933	2+2-	INS	-108	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19350782	2+0-	20	19350974	0+3-	INS	-140	19	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	19356433	3+2-	20	19356456	3+2-	INS	-207	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19357097	2+2-	20	19357111	2+2-	INS	-209	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19366367	2+0-	20	19366360	0+2-	INS	-342	27	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	19370055	2+2-	20	19370076	2+2-	INS	-213	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19388317	2+2-	20	19388338	2+2-	INS	-228	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19395628	2+0-	20	19395704	3+5-	INS	-143	38	4	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19419731	3+0-	20	19419813	1+5-	INS	-172	35	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	19423485	2+2-	20	19423461	2+2-	INS	-391	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19427244	2+2-	20	19427265	2+2-	INS	-92	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19430347	2+2-	20	19430390	0+2-	INS	-247	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19438548	2+3-	20	19438559	2+3-	INS	-230	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19439690	3+1-	20	19439801	2+3-	INS	-207	29	3	COLO-829_v2_74|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	19447001	2+2-	20	19446996	2+2-	INS	-88	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19455314	2+0-	20	19455406	0+2-	INS	-223	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19467212	2+3-	20	19467262	2+3-	INS	-194	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19472067	3+1-	20	19472218	0+2-	INS	-128	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19487399	2+2-	20	19487418	2+2-	INS	-95	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19489954	3+0-	20	19490012	0+2-	INS	-267	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19490982	4+4-	20	19491027	4+4-	INS	-100	53	4	COLO-829-IL|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19500052	2+0-	20	19500095	0+2-	INS	-268	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19503124	3+4-	20	19503153	3+4-	INS	-183	29	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19507418	2+2-	20	19507463	2+2-	INS	-95	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19507985	2+2-	20	19507985	2+2-	INS	-97	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19520225	2+2-	20	19520238	2+2-	INS	-382	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19528478	3+3-	20	19528461	3+3-	INS	-366	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19528694	2+3-	20	19528699	2+3-	INS	-109	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19533688	3+4-	20	19533808	3+4-	INS	-212	19	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19540344	2+4-	20	19540331	2+4-	INS	-97	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19558341	2+0-	20	19558346	0+2-	INS	-200	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	19569793	3+1-	20	19569871	1+5-	INS	-217	37	4	COLO-829_v2_74|4	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	19582605	2+3-	20	19582593	2+3-	INS	-103	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19589280	2+2-	20	19589296	2+2-	INS	-209	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19595638	2+2-	20	19595665	2+2-	INS	-103	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19599335	2+0-	20	19599416	0+2-	INS	-241	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19609386	3+2-	20	19609419	3+2-	INS	-341	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19610148	2+3-	20	19610219	2+3-	INS	-217	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19612510	3+1-	20	19612626	0+3-	INS	-140	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	19618408	3+2-	20	19618480	3+2-	INS	-92	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19676293	3+2-	20	19676318	3+2-	INS	-103	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19691753	2+2-	20	19691741	2+2-	INS	-107	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	19698643	2+2-	20	19698695	2+2-	INS	-88	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19703451	2+2-	20	19703417	2+2-	INS	-109	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19732714	2+2-	20	19732676	2+2-	INS	-108	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19736215	2+1-	20	19736367	0+2-	INS	-151	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19737493	2+2-	20	19737488	2+2-	INS	-245	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19746919	2+3-	20	19746982	2+3-	INS	-321	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19751509	14+13-	20	19754808	1+16-	DEL	3305	99	14	COLO-829BL-IL|2:COLO-829-IL|12	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	19751509	0+13-	20	19754262	4+2-	ITX	2393	83	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19751509	0+10-	20	19754560	9+1-	ITX	2906	99	9	COLO-829BL-IL|4:COLO-829-IL|5	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	19773274	4+8-	20	19773314	4+8-	INS	-88	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	19779722	11+0-	20	19779722	0+2-	INS	-182	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19786033	3+2-	20	19786057	3+2-	INS	-99	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19790020	2+2-	20	19789981	2+2-	INS	-388	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19793470	2+2-	20	19793476	2+2-	INS	-219	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19800736	2+2-	20	19800700	2+2-	INS	-249	26	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19804366	2+0-	20	19804489	1+2-	INS	-164	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19845293	2+0-	20	19845355	0+2-	INS	-250	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19853028	3+2-	20	19853067	12+14-	INS	-295	99	11	COLO-829_v2_74|9:COLO-829-IL|2	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	19862989	3+4-	20	19863016	3+4-	INS	-375	28	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19866079	2+2-	20	19866100	2+2-	INS	-100	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19918396	2+1-	20	19918524	0+2-	INS	-161	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19930412	2+2-	20	19930393	2+2-	INS	-88	33	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19944139	2+2-	20	19944119	2+2-	INS	-370	22	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	19950484	2+1-	20	19950587	0+2-	INS	-161	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	19960256	3+0-	20	19960388	0+2-	INS	-163	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19971560	2+0-	20	19971651	1+2-	INS	-249	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20009791	2+2-	20	20009804	2+2-	INS	-99	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20013798	3+0-	20	20014003	0+2-	INS	-114	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20016399	2+2-	20	20016391	2+2-	INS	-235	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20022665	3+2-	20	20022706	0+2-	INS	-252	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20033873	2+2-	20	20033850	2+2-	INS	-401	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20034197	2+2-	20	20034179	2+2-	INS	-91	29	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20035133	2+2-	20	20035144	2+2-	INS	-101	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20046128	2+3-	20	20046126	2+3-	INS	-122	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20062359	2+0-	20	20062462	0+3-	INS	-215	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	19463041	13+0-	20	20104120	30+32-	DEL	641076	80	4	COLO-829BL-IL|2:COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	19463234	1+9-	20	20104120	29+27-	ITX	640706	76	4	COLO-829BL-IL|1:COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20086077	2+2-	20	20086076	2+2-	INS	-94	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20111924	2+2-	20	20111883	2+2-	INS	-390	27	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20114029	2+3-	20	20114041	2+3-	INS	-113	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20135272	3+3-	20	20135246	3+3-	INS	-376	38	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20145979	2+2-	20	20145945	2+2-	INS	-107	32	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20159917	2+1-	20	20160051	0+2-	INS	-183	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20167788	2+2-	20	20167767	2+2-	INS	-371	22	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20174246	3+1-	20	20174243	1+2-	INS	-198	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20177609	2+2-	20	20177657	2+2-	INS	-235	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20178785	2+2-	20	20178820	2+2-	INS	-242	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20182317	2+3-	20	20182376	2+3-	INS	-337	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20182785	2+0-	20	20182900	0+2-	DEL	93	40	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20184151	2+2-	20	20184140	2+2-	ITX	-129	41	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20219321	2+1-	20	20219326	1+3-	INS	-143	28	3	COLO-829_v2_74|1:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20224567	15+11-	20	20224917	15+11-	DEL	90	99	7	COLO-829BL-IL|5:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	20226629	2+2-	20	20226630	2+2-	INS	-227	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20235742	4+3-	20	20235791	4+3-	INS	-108	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20246150	2+4-	20	20246173	2+4-	INS	-109	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20249109	2+0-	20	20249245	1+3-	DEL	92	41	2	COLO-829-IL|2	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	20260150	2+1-	20	20260182	1+3-	INS	-334	24	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	20265820	306+287-	20	20266228	306+287-	ITX	-153	99	111	COLO-829BL-IL|45:COLO-829_v2_74|1:COLO-829-IL|65	0.27	BreakDancerMax-0.0.1r81	|q10|o20
20	20266298	56+37-	20	20266283	1+36-	DEL	141	99	33	COLO-829BL-IL|12:COLO-829-IL|21	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	20283976	3+0-	20	20284010	16+20-	INS	-293	65	9	COLO-829BL-IL|1:COLO-829_v2_74|6:COLO-829-IL|2	0.60	BreakDancerMax-0.0.1r81	|q10|o20
20	20284321	6+8-	20	20284995	46+39-	ITX	-84	99	24	COLO-829BL-IL|12:COLO-829-IL|12	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	20284321	5+5-	20	20284456	3+3-	ITX	-29	44	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20284321	4+2-	20	20286406	18+23-	ITX	233	99	10	COLO-829BL-IL|4:COLO-829_v2_74|3:COLO-829-IL|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	20285234	15+10-	20	20286406	8+14-	DEL	1362	99	11	COLO-829BL-IL|1:COLO-829-IL|10	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	20285234	4+2-	20	20285236	0+2-	DEL	92	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	20285234	2+2-	20	20285709	2+3-	DEL	468	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	20285832	2+1-	20	20286406	0+3-	DEL	392	39	2	COLO-829_v2_74|2	0.29	BreakDancerMax-0.0.1r81	|q10|o20
20	20284951	1+9-	20	20285587	12+5-	ITX	330	99	11	COLO-829BL-IL|7:COLO-829-IL|4	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	20311921	2+1-	20	20311986	1+2-	INS	-252	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20327543	2+2-	20	20327556	2+2-	INS	-108	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20355014	2+2-	20	20355013	2+2-	INS	-104	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20370674	2+0-	20	20370671	0+2-	INS	-329	23	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20378044	3+3-	20	20378091	3+3-	INS	-112	22	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20429272	4+0-	20	20429263	1+2-	INS	-326	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20442712	2+2-	20	20442699	2+2-	INS	-118	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20442946	2+2-	20	20442988	2+2-	INS	-198	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20450723	2+3-	20	20450745	2+3-	INS	-111	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20456942	2+2-	20	20456891	2+2-	INS	-122	38	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20477562	2+2-	20	20477620	2+2-	INS	-212	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20485532	2+2-	20	20485484	2+2-	INS	-398	29	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20490137	2+2-	20	20490124	2+2-	INS	-118	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20495260	3+3-	20	20495275	3+3-	INS	-95	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20497533	2+0-	20	20497533	1+3-	INS	-207	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	20512232	2+2-	20	20512239	2+2-	INS	-223	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20515157	2+0-	20	20515278	0+2-	INS	-198	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20520437	2+3-	20	20520470	2+3-	INS	-245	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20535740	2+2-	20	20535703	2+2-	INS	-386	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20535927	3+1-	20	20536008	0+2-	INS	-248	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20545857	2+0-	20	20546002	1+3-	INS	-161	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20551637	4+2-	20	20551611	4+2-	INS	-121	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20567741	2+2-	20	20567726	2+2-	INS	-110	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20570484	3+1-	20	20570624	0+2-	INS	-136	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20583645	2+2-	20	20583662	2+2-	INS	-97	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20598733	2+3-	20	20598808	2+3-	INS	-233	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20610545	2+2-	20	20610551	2+2-	INS	-255	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20615042	2+2-	20	20615002	2+2-	INS	-114	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20615501	2+3-	20	20615532	2+3-	INS	-228	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20618902	2+0-	20	20619036	0+2-	INS	-186	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20627715	2+2-	20	20627720	2+2-	INS	-95	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20656084	3+1-	20	20656221	0+2-	INS	-146	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20660375	2+0-	20	20660508	0+2-	INS	-178	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20677990	2+0-	20	20678058	4+7-	INS	-136	33	6	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	20679445	2+2-	20	20679414	2+2-	INS	-380	24	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20691242	3+2-	20	20691275	3+2-	INS	-115	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20700000	2+1-	20	20700068	0+2-	INS	-229	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20715709	2+0-	20	20715766	1+4-	INS	-191	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20749053	3+1-	20	20749116	0+4-	INS	-224	23	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20754873	5+5-	20	20754976	5+5-	INS	-154	36	4	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20756635	7+1-	20	20756643	0+8-	DEL	88	99	6	COLO-829BL-IL|2:COLO-829-IL|4	0.17	BreakDancerMax-0.0.1r81	|q10|o20
20	20770864	2+2-	20	20770814	2+2-	INS	-116	41	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20785427	2+2-	20	20785442	2+2-	INS	-104	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20785943	2+3-	20	20785978	2+3-	INS	-100	27	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20792024	3+2-	20	20792203	3+2-	INS	-122	24	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20792336	3+0-	20	20792459	0+4-	INS	-225	30	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20805894	4+2-	20	20805927	4+2-	INS	-208	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20808942	2+3-	20	20808924	2+3-	INS	-106	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20809198	2+0-	20	20809364	0+3-	INS	-149	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20812513	4+2-	20	20812556	4+2-	INS	-103	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20812626	2+0-	20	20812654	0+2-	INS	-212	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20818698	2+2-	20	20818680	2+2-	INS	-100	33	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20820612	2+0-	20	20820667	0+2-	INS	-275	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20830749	2+2-	20	20830716	2+2-	INS	-102	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	20845844	2+2-	20	20845801	2+2-	INS	-393	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20849453	2+1-	20	20849686	1+2-	INS	-106	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20849946	2+0-	20	20849976	0+3-	INS	-274	16	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20855395	2+0-	20	20855572	0+2-	INS	-142	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20882707	3+1-	20	20882818	0+2-	INS	-171	39	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20890367	6+1-	20	20890397	1+7-	INS	-216	60	7	COLO-829_v2_74|6:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	20904247	3+1-	20	20904384	0+2-	INS	-272	44	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20910410	2+3-	20	20910391	2+3-	INS	-392	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20911009	2+2-	20	20910969	2+2-	INS	-103	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20943966	3+5-	20	20944141	3+5-	INS	-162	10	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20952466	2+1-	20	20952484	1+2-	INS	-292	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20956690	4+2-	20	20956774	4+2-	INS	-92	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20958159	3+0-	20	20958243	0+3-	INS	-236	30	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	20958727	2+0-	20	20958913	0+2-	INS	-146	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	20970213	2+2-	20	20970201	2+2-	INS	-99	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	20978761	2+1-	20	20978763	1+3-	INS	-248	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	21013324	2+0-	20	21013413	0+2-	INS	-218	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21018336	3+4-	20	21018380	3+4-	INS	-272	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21024644	2+2-	20	21024655	2+2-	INS	-87	29	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21041127	2+2-	20	21041146	2+2-	INS	-105	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21047560	2+2-	20	21047575	2+2-	INS	-98	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21050503	2+6-	20	21050645	2+6-	INS	-304	11	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21072227	2+0-	20	21072414	0+2-	INS	-140	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21077504	3+3-	20	21077559	3+3-	INS	-184	26	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21079663	2+2-	20	21079662	2+2-	INS	-99	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21080757	2+1-	20	21080808	0+2-	INS	-235	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21089880	4+3-	20	21089925	1+2-	INS	-201	29	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21091746	2+3-	20	21091779	2+3-	INS	-230	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21102722	2+3-	20	21102770	2+3-	INS	-95	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21122794	2+2-	20	21122739	2+2-	INS	-117	38	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21151303	2+2-	20	21151306	2+2-	INS	-222	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21201945	3+3-	20	21201985	3+3-	INS	-364	27	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21214992	2+0-	20	21215044	0+2-	INS	-281	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21216505	2+5-	20	21216484	2+5-	INS	-113	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21222579	2+0-	20	21222613	1+3-	INS	-242	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	21228389	3+0-	20	21228475	0+3-	INS	-253	48	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21233828	5+0-	20	21236755	2+67-	DEL	2693	86	4	COLO-829_v2_74|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	21234133	66+0-	20	21236755	0+61-	DEL	2680	99	61	COLO-829BL-IL|23:COLO-829_v2_74|3:COLO-829-IL|35	0.61	BreakDancerMax-0.0.1r81	|q10|o20
20	21244420	3+2-	20	21244467	3+2-	INS	-243	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21247375	2+2-	20	21247340	2+2-	INS	-243	25	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21264043	2+2-	20	21264006	2+2-	INS	-100	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21276155	2+2-	20	21276166	2+2-	INS	-227	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21291517	2+2-	20	21291521	2+2-	INS	-103	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21301628	3+3-	20	21301629	3+3-	INS	-101	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21314127	2+3-	20	21314178	2+3-	INS	-208	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21315508	2+2-	20	21315474	2+2-	INS	-106	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21330701	2+2-	20	21330653	2+2-	INS	-119	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21340759	2+2-	20	21340741	2+2-	INS	-109	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21350372	2+2-	20	21350366	2+2-	INS	-98	27	2	COLO-829-IL|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	21353483	2+0-	20	21353588	1+3-	INS	-180	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	21365994	2+2-	20	21366002	2+2-	INS	-373	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21377524	4+4-	20	21377651	4+4-	INS	-98	17	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21380502	3+2-	20	21380527	3+2-	INS	-247	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21383758	2+2-	20	21383764	2+2-	INS	-226	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21385080	2+2-	20	21385088	2+2-	INS	-98	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21395437	2+0-	20	21395509	0+2-	INS	-252	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21395873	2+3-	20	21395907	2+3-	INS	-111	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21412471	2+2-	20	21412508	2+2-	INS	-109	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21417338	2+2-	20	21417309	2+2-	INS	-106	35	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21453364	2+2-	20	21453373	2+2-	INS	-252	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21465465	3+2-	20	21465470	0+2-	INS	-181	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21468754	2+2-	20	21468712	2+2-	INS	-115	34	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21472880	3+0-	20	21472978	1+3-	INS	-189	45	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21484030	2+2-	20	21483993	2+2-	INS	-387	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21488829	2+3-	20	21488831	2+3-	INS	-218	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21512359	2+2-	20	21512353	2+2-	INS	-230	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21512553	3+2-	20	21512615	3+2-	INS	-343	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21514342	3+0-	20	21514371	1+4-	INS	-229	43	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	21520021	2+2-	20	21520018	2+2-	INS	-113	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21529637	2+2-	20	21529595	2+2-	INS	-119	34	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21530699	2+2-	20	21530680	2+2-	INS	-105	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21591588	2+3-	20	21591628	2+3-	INS	-228	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21597691	2+2-	20	21597731	2+2-	INS	-92	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21607791	2+3-	20	21607881	2+3-	INS	-253	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21613114	2+3-	20	21613108	2+3-	INS	-90	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21624173	2+1-	20	21624257	0+2-	INS	-241	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21641313	2+3-	20	21641293	2+3-	INS	-102	33	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21650276	23+23-	20	21650317	23+23-	INS	-106	99	14	COLO-829BL-IL|6:COLO-829-IL|8	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21664720	2+0-	20	21664861	0+2-	INS	-167	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21669804	3+1-	20	21669871	0+3-	INS	-154	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21707297	2+2-	20	21707324	2+2-	INS	-248	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21708523	2+0-	20	21708619	0+3-	INS	-197	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21710690	2+2-	20	21710682	2+2-	INS	-109	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21712397	2+1-	20	21712435	1+2-	INS	-261	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21729866	2+0-	20	21729930	3+4-	INS	-167	34	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21741175	2+0-	20	21741211	1+3-	INS	-199	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	21752015	2+2-	20	21752015	2+2-	INS	-384	19	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21772919	2+2-	20	21772899	2+2-	INS	-244	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21775518	2+2-	20	21775523	2+2-	INS	-94	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21777943	3+1-	20	21777992	1+2-	INS	-222	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	21793570	2+2-	20	21793543	2+2-	INS	-93	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21794858	2+2-	20	21794846	2+2-	INS	-91	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21797630	5+0-	20	21798184	0+60-	DEL	282	99	5	COLO-829_v2_74|5	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	21797955	66+3-	20	21798184	0+55-	DEL	291	99	55	COLO-829BL-IL|16:COLO-829-IL|39	0.53	BreakDancerMax-0.0.1r81	|q10|o20
20	21797955	8+0-	20	21798425	1+7-	DEL	294	99	7	COLO-829_v2_74|7	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	21819424	10+0-	20	21842263	23+18-	INV	22748	99	10	COLO-829BL-IL|5:COLO-829-IL|5	0.62	BreakDancerMax-0.0.1r81	|q10|o20
20	21822310	4+6-	20	21822308	0+3-	INS	-87	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	21823759	2+2-	20	21823728	2+2-	INS	-113	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	21832487	3+0-	20	21832543	0+2-	INS	-248	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21848496	2+2-	20	21848509	2+2-	INS	-233	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21860395	8+14-	20	21860527	8+14-	INS	-110	17	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	21879872	3+3-	20	21879865	3+3-	INS	-111	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21880966	2+3-	20	21880956	2+3-	INS	-104	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21891539	2+0-	20	21891736	0+2-	INS	-115	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21892428	2+3-	20	21892423	2+3-	INS	-121	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21897387	3+2-	20	21897413	0+3-	INS	-304	29	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21905210	3+3-	20	21905249	3+3-	INS	-232	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21910693	2+0-	20	21910724	0+2-	INS	-290	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21941557	5+2-	20	21941571	5+2-	INS	-105	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	21946565	2+2-	20	21946547	2+2-	INS	-254	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21960924	2+2-	20	21960888	2+2-	INS	-101	33	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21963868	2+2-	20	21963846	2+2-	INS	-252	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	21977705	14+15-	20	21977804	14+15-	INS	-95	19	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	21987145	3+2-	20	21987132	3+2-	INS	-227	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21996982	2+2-	20	21996940	2+2-	INS	-108	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	21997672	3+3-	20	21997669	3+3-	INS	-286	34	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	21999350	3+2-	20	21999363	3+2-	INS	-212	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22002011	2+2-	20	22001989	2+2-	INS	-102	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22020355	3+1-	20	22020489	0+2-	INS	-164	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22042685	2+2-	20	22042635	2+2-	INS	-119	37	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22065409	2+2-	20	22065417	2+2-	INS	-99	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22076858	3+4-	20	22076889	3+4-	INS	-252	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22082166	2+2-	20	22082167	2+2-	INS	-229	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	22089142	2+2-	20	22089168	2+2-	INS	-99	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22102726	2+2-	20	22102694	2+2-	INS	-104	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22106710	2+2-	20	22106727	2+2-	INS	-106	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22107063	3+1-	20	22107112	2+4-	INS	-159	43	5	COLO-829_v2_74|2:COLO-829-IL|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	22122141	2+2-	20	22122094	2+2-	INS	-119	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22155718	2+0-	20	22155782	0+3-	INS	-258	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22182277	2+2-	20	22182263	2+2-	INS	-253	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22188660	2+5-	20	22188653	2+5-	ITX	-126	41	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22194515	2+2-	20	22194506	2+2-	INS	-240	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	22203265	3+2-	20	22203289	3+2-	INS	-105	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22217638	3+1-	20	22217717	0+2-	INS	-250	25	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22239675	2+2-	20	22239648	2+2-	INS	-95	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22239868	2+1-	20	22239864	0+2-	INS	-311	18	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	22253952	3+0-	20	22254067	1+3-	INS	-229	38	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22264226	2+2-	20	22264259	2+2-	INS	-91	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22286744	2+0-	20	22286734	0+2-	INS	-336	23	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	22297485	3+4-	20	22297585	3+4-	INS	-259	22	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22340032	2+2-	20	22340012	2+2-	INS	-110	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	22359848	2+2-	20	22359827	2+2-	INS	-371	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22362966	2+2-	20	22362938	2+2-	INS	-99	35	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22364073	3+3-	20	22364127	3+3-	INS	-166	28	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22377761	2+2-	20	22377797	2+2-	INS	-221	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22383383	2+2-	20	22383353	2+2-	INS	-95	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	22384451	2+2-	20	22384541	0+2-	INS	-241	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22395012	2+3-	20	22395072	2+3-	INS	-371	15	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	22400593	2+0-	20	22400580	0+2-	INS	-91	32	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	22412365	2+2-	20	22412334	2+2-	INS	-102	36	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22414438	2+3-	20	22414457	2+3-	INS	-109	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22429843	2+0-	20	22430056	0+2-	INS	-124	28	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22434161	27+2-	20	22434183	10+14-	DEL	97	99	10	COLO-829BL-IL|4:COLO-829-IL|6	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	22454561	2+3-	20	22454676	0+2-	INS	-210	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22455509	2+2-	20	22455453	2+2-	INS	-406	33	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	22456795	10+2-	20	22456851	10+2-	INS	-113	22	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	22467292	2+0-	20	22467603	0+19-	DEL	104	46	2	COLO-829_v2_74|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	22467522	22+1-	20	22467603	0+17-	DEL	95	99	13	COLO-829BL-IL|3:COLO-829-IL|10	0.45	BreakDancerMax-0.0.1r81	|q10|o20
20	22467522	9+1-	20	22467834	0+5-	DEL	87	99	5	COLO-829_v2_74|5	0.24	BreakDancerMax-0.0.1r81	|q10|o20
20	22475220	3+0-	20	22475214	1+3-	INS	-281	26	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	22483123	3+1-	20	22483183	0+2-	INS	-208	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22501796	2+2-	20	22501779	2+2-	INS	-102	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22517335	2+0-	20	22517411	2+5-	INS	-139	20	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	22520809	3+2-	20	22520872	3+2-	INS	-97	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22529433	2+2-	20	22529412	2+2-	INS	-109	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22530281	3+2-	20	22530297	3+2-	INS	-100	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22534613	3+4-	20	22534629	3+4-	INS	-286	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22543487	2+2-	20	22543459	2+2-	INS	-90	35	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22547123	2+0-	20	22547131	1+3-	INS	-215	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	22548015	2+0-	20	22548103	0+2-	INS	-239	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22565734	2+2-	20	22565748	2+2-	INS	-103	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22566246	2+2-	20	22566214	2+2-	INS	-108	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22571365	3+3-	20	22571436	3+3-	INS	-193	25	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22602086	4+1-	20	22602137	1+5-	INS	-221	38	5	COLO-829_v2_74|5	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22603364	36+0-	20	22604006	0+2-	DEL	345	44	2	COLO-829_v2_74|2	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	22603364	34+0-	20	22603648	0+34-	DEL	340	99	32	COLO-829BL-IL|14:COLO-829-IL|18	0.63	BreakDancerMax-0.0.1r81	|q10|o20
20	22633880	3+4-	20	22633914	3+4-	INS	-120	35	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22638983	2+2-	20	22638935	2+2-	INS	-397	29	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	22639522	2+0-	20	22639565	1+3-	INS	-202	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22656595	2+2-	20	22656609	2+2-	INS	-93	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22659120	2+2-	20	22659139	2+2-	INS	-221	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22676893	2+2-	20	22676882	2+2-	INS	-110	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22700566	2+3-	20	22700563	2+3-	INS	-106	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	22707741	2+3-	20	22707822	2+3-	INS	-183	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22715229	2+4-	20	22715265	2+4-	INS	-325	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22719493	2+2-	20	22719493	2+2-	INS	-114	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22724383	2+3-	20	22724375	2+3-	INS	-110	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	22747586	2+3-	20	22747636	2+3-	INS	-87	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22754826	3+2-	20	22754905	3+2-	INS	-88	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22755374	2+0-	20	22755412	0+3-	INS	-258	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22773196	2+2-	20	22773227	2+2-	INS	-98	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22782997	2+3-	20	22783041	2+3-	INS	-100	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22789739	3+0-	20	22789815	0+2-	INS	-231	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22790614	2+2-	20	22790597	2+2-	INS	-102	33	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22795860	2+2-	20	22795815	2+2-	INS	-116	35	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22808972	3+1-	20	22809126	0+3-	INS	-162	31	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22811387	6+10-	20	22811553	6+10-	INS	-91	54	5	COLO-829-IL|5	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	22813069	2+2-	20	22813087	2+2-	INS	-95	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22820442	3+2-	20	22820448	3+2-	INS	-253	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22834193	3+0-	20	22834288	0+3-	INS	-235	35	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22842769	3+2-	20	22842754	3+2-	INS	-101	33	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22874092	2+0-	20	22874195	0+2-	INS	-246	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22876977	2+2-	20	22877020	2+2-	INS	-194	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22889430	3+3-	20	22889437	3+3-	INS	-228	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22890045	2+0-	20	22890176	0+2-	INS	-145	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22893574	2+6-	20	22893658	2+6-	INS	-195	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22901695	3+2-	20	22901692	3+2-	INS	-96	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22902787	2+2-	20	22902796	2+2-	INS	-227	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22908028	3+2-	20	22908036	3+2-	INS	-107	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22928558	2+2-	20	22928528	2+2-	INS	-105	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22933471	2+3-	20	22933505	2+3-	INS	-98	23	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	22959378	2+1-	20	22959401	0+3-	INS	-258	14	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22972362	2+2-	20	22972365	2+2-	INS	-100	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22981939	3+2-	20	22981974	3+2-	INS	-93	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	22989665	2+3-	20	22989678	2+3-	INS	-107	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22992751	2+3-	20	22992718	2+3-	INS	-118	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	22993409	2+2-	20	22993389	2+2-	INS	-102	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	22998354	2+2-	20	22998317	2+2-	INS	-100	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	23008614	2+2-	20	23008592	2+2-	INS	-105	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23022527	2+2-	20	23022488	2+2-	INS	-389	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23025959	2+0-	20	23026134	0+2-	INS	-145	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23028077	3+1-	20	23028181	0+2-	INS	-176	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23033466	2+2-	20	23033452	2+2-	INS	-94	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23035004	2+2-	20	23035007	2+2-	INS	-255	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23051301	25+2-	20	23051633	0+14-	DEL	299	99	14	COLO-829BL-IL|2:COLO-829_v2_74|8:COLO-829-IL|4	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	23051301	8+1-	20	23051804	0+8-	DEL	310	99	8	COLO-829_v2_74|8	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	23053362	2+0-	20	23053465	1+3-	INS	-173	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23064777	2+3-	20	23064807	2+3-	INS	-106	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23073343	2+0-	20	23073486	0+2-	INS	-165	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23076621	3+3-	20	23076630	3+3-	INS	-207	33	3	COLO-829_v2_74|1:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	23080352	3+1-	20	23080543	1+3-	INS	-108	39	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23081017	2+2-	20	23080958	2+2-	INS	-409	35	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23084329	4+2-	20	23084434	2+3-	INS	-94	23	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23096149	2+0-	20	23096234	0+2-	INS	-222	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23133898	2+0-	20	23133918	0+2-	INS	-260	18	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	23159423	3+3-	20	23159447	3+3-	INS	-101	37	3	COLO-829BL-IL|1:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23160058	2+2-	20	23160085	2+2-	INS	-206	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23161242	2+2-	20	23161230	2+2-	INS	-241	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23176965	2+3-	20	23176999	2+3-	INS	-241	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23203964	2+0-	20	23204151	0+2-	INS	-142	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23214947	2+2-	20	23214951	2+2-	INS	-236	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23218946	2+3-	20	23218978	2+3-	INS	-366	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23237617	2+2-	20	23237612	2+2-	INS	-100	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23242112	2+1-	20	23242256	0+2-	INS	-152	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23243334	33+33-	20	23243396	33+33-	INS	-103	99	29	COLO-829BL-IL|14:COLO-829-IL|15	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	23250813	3+1-	20	23250983	0+2-	INS	-205	27	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23254047	2+3-	20	23254101	2+3-	INS	-249	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23272943	2+3-	20	23272917	2+3-	INS	-100	31	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23278642	2+2-	20	23278604	2+2-	INS	-107	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23282328	2+0-	20	23282468	0+3-	INS	-194	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23288197	2+2-	20	23288179	2+2-	INS	-101	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23288574	2+2-	20	23288554	2+2-	INS	-118	33	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23292210	3+2-	20	23292247	3+2-	INS	-347	16	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	23301498	2+3-	20	23301523	2+3-	INS	-219	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23305966	3+4-	20	23306102	3+4-	INS	-198	22	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23306558	2+3-	20	23306535	2+3-	INS	-99	34	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23319664	2+2-	20	23319644	2+2-	INS	-96	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23365371	2+2-	20	23365386	2+2-	INS	-89	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23380816	2+3-	20	23380827	2+3-	INS	-257	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	23388410	2+1-	20	23388489	1+2-	INS	-270	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23416864	3+3-	20	23416899	3+3-	INS	-100	37	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23429157	3+1-	20	23429212	1+3-	INS	-265	41	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	23433455	3+0-	20	23433560	5+3-	INS	-153	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	23450443	2+5-	20	23450529	2+5-	INS	-227	15	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23477639	2+3-	20	23477632	2+3-	INS	-254	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	23489359	2+0-	20	23489743	1+16-	DEL	101	47	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23489719	23+13-	20	23489743	0+13-	DEL	97	99	11	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|8	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	23494064	2+0-	20	23494121	0+2-	INS	-277	27	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23495138	2+2-	20	23495098	2+2-	INS	-104	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23498273	3+2-	20	23498287	3+2-	INS	-234	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23499193	2+3-	20	23499207	2+3-	INS	-258	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23502562	8+3-	20	23502569	8+3-	INS	-266	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	23505126	2+2-	20	23505110	2+2-	INS	-91	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23512568	2+2-	20	23512585	2+2-	INS	-102	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23516121	2+2-	20	23516083	2+2-	INS	-249	26	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23558102	3+3-	20	23558091	3+3-	INS	-97	44	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23565542	2+2-	20	23565510	2+2-	INS	-244	27	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23572934	3+0-	20	23573019	0+2-	INS	-218	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23582125	3+2-	20	23582167	3+2-	INS	-93	27	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	23588833	2+1-	20	23588892	0+3-	INS	-231	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23589882	2+1-	20	23589975	0+2-	INS	-209	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23595068	2+2-	20	23595044	2+2-	INS	-374	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23604973	2+3-	20	23604992	2+3-	INS	-233	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23606280	3+0-	20	23661556	0+3-	DEL	55268	56	3	COLO-829BL-IL|1:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	23613843	2+1-	20	23675755	0+2-	DEL	61751	41	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23620776	2+2-	20	23620731	2+2-	INS	-395	28	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23664177	3+3-	20	23664208	3+3-	INS	-111	39	3	COLO-829-IL|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23630788	4+6-	20	23774893	0+3-	DEL	144077	58	3	COLO-829BL-IL|1:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23630788	1+6-	20	23774608	6+1-	ITX	143650	99	6	COLO-829BL-IL|3:COLO-829-IL|3	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	23655796	5+1-	20	23731531	18+3-	DEL	75774	52	3	COLO-829BL-IL|1:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23656005	0+19-	20	23731531	18+0-	ITX	75407	99	18	COLO-829BL-IL|6:COLO-829-IL|12	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	23662692	4+0-	20	23738476	14+4-	DEL	75817	82	4	COLO-829BL-IL|3:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	23662909	1+13-	20	23738476	14+0-	ITX	75427	99	13	COLO-829BL-IL|3:COLO-829-IL|10	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	23667637	8+0-	20	23743548	11+8-	DEL	75885	99	8	COLO-829BL-IL|2:COLO-829-IL|6	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	23667901	0+11-	20	23743548	11+0-	ITX	75487	99	11	COLO-829BL-IL|6:COLO-829-IL|5	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23677482	4+1-	20	23753685	4+4-	DEL	76189	79	4	COLO-829BL-IL|1:COLO-829-IL|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	23677689	0+3-	20	23753685	4+0-	ITX	75814	67	3	COLO-829BL-IL|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23701249	2+0-	20	23701398	0+2-	INS	-160	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23702840	3+0-	20	23702917	0+2-	INS	-234	19	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23735952	4+2-	20	23736039	4+2-	INS	-100	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23749420	5+3-	20	23749494	5+3-	INS	-112	34	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23749564	2+0-	20	23749552	1+3-	INS	-162	21	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23752439	2+2-	20	23752417	2+2-	INS	-103	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23755305	3+4-	20	23755323	3+4-	INS	-116	37	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23766652	2+2-	20	23766646	2+2-	INS	-98	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23775072	2+2-	20	23775054	2+2-	INS	-243	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23705136	0+2-	20	23786602	2+0-	ITX	81288	42	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23781109	2+2-	20	23781088	2+2-	INS	-110	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23806448	4+3-	20	23806483	4+3-	INS	-213	34	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23817907	3+2-	20	23817917	3+2-	INS	-116	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	23822063	2+2-	20	23822025	2+2-	INS	-387	26	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23829357	3+4-	20	23829338	3+4-	INS	-103	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	23833059	2+0-	20	23833232	1+4-	INS	-120	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23834503	3+3-	20	23834537	3+3-	INS	-275	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23834808	2+0-	20	23834921	0+2-	INS	-202	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23842385	2+0-	20	23842561	0+2-	INS	-141	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23845248	3+4-	20	23845254	3+4-	INS	-353	31	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23848367	3+3-	20	23848461	3+3-	INS	-378	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23843109	2+0-	20	23883110	14+11-	DEL	39712	51	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	23843396	9+1-	20	23883110	14+9-	DEL	39724	99	9	COLO-829BL-IL|3:COLO-829-IL|6	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	23843639	0+13-	20	23883110	14+0-	ITX	39330	99	13	COLO-829BL-IL|6:COLO-829-IL|7	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	23871300	19+3-	20	23871283	2+20-	INS	-146	99	17	COLO-829BL-IL|1:COLO-829_v2_74|13:COLO-829-IL|3	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	23886316	2+2-	20	23886257	2+2-	INS	-409	35	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23900514	2+2-	20	23900532	2+2-	INS	-100	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23959179	2+0-	20	23959246	0+2-	INS	-253	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23963807	2+0-	20	23963873	0+2-	INS	-246	19	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	23966223	2+1-	20	23966280	1+3-	INS	-209	34	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23971987	3+1-	20	23972030	0+2-	INS	-203	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23975283	3+3-	20	23975357	3+3-	INS	-105	34	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23982892	2+1-	20	23982979	0+2-	INS	-223	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	23989909	3+0-	20	23990011	0+3-	INS	-230	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	23995720	2+4-	20	23995792	2+4-	INS	-102	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24009744	2+2-	20	24009708	2+2-	INS	-386	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24027536	2+3-	20	24027609	2+3-	INS	-92	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24029210	2+2-	20	24029190	2+2-	INS	-251	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24067872	2+2-	20	24067851	2+2-	INS	-371	22	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24069543	2+2-	20	24069507	2+2-	INS	-122	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24077022	3+0-	20	24077110	0+2-	INS	-240	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24079289	2+2-	20	24079247	2+2-	INS	-112	34	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24081382	2+2-	20	24081363	2+2-	INS	-254	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24103708	2+2-	20	24103676	2+2-	INS	-99	36	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24110937	2+3-	20	24110935	2+3-	INS	-99	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24122249	3+1-	20	24122329	1+3-	INS	-209	23	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24127038	4+3-	20	24127131	4+3-	INS	-105	30	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24134804	2+2-	20	24134773	2+2-	INS	-255	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24136547	3+0-	20	24137035	1+5-	DEL	231	70	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	24138708	2+0-	20	24138856	0+2-	INS	-158	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24160924	3+1-	20	24161028	2+4-	INS	-165	58	5	COLO-829_v2_74|2:COLO-829-IL|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	24163957	3+1-	20	24164103	0+2-	INS	-247	29	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24169056	3+3-	20	24169074	3+3-	INS	-120	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24190951	3+3-	20	24190957	3+3-	INS	-92	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24229521	2+2-	20	24229537	2+2-	INS	-240	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24230867	2+2-	20	24230828	2+2-	INS	-388	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24235809	2+2-	20	24235824	2+2-	INS	-115	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24262680	2+2-	20	24262625	2+2-	INS	-405	32	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24275565	3+3-	20	24275530	3+3-	INS	-104	51	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24285634	3+3-	20	24285636	3+3-	INS	-102	43	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24303728	3+3-	20	24303758	3+3-	INS	-290	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24305443	2+2-	20	24305456	2+2-	INS	-103	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24308603	2+2-	20	24308634	2+2-	INS	-90	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24325693	2+4-	20	24325726	2+4-	INS	-123	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24337477	2+0-	20	24337539	2+3-	DEL	91	42	2	COLO-829BL-IL|2	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	24347740	2+2-	20	24347722	2+2-	INS	-105	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24360034	3+1-	20	24360153	0+4-	DEL	90	51	3	COLO-829BL-IL|1:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	24386214	3+3-	20	24386290	3+3-	INS	-93	31	3	COLO-829BL-IL|1:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24416066	2+0-	20	24416225	0+2-	INS	-163	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24421015	2+2-	20	24420992	2+2-	INS	-98	34	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24433814	2+2-	20	24433839	2+2-	INS	-89	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24441783	2+3-	20	24441774	2+3-	INS	-101	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24458574	28+27-	20	24458732	28+27-	INS	-92	99	21	COLO-829BL-IL|7:COLO-829-IL|14	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	24464878	2+2-	20	24464846	2+2-	INS	-394	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24497231	2+2-	20	24497259	2+2-	INS	-249	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24505830	2+1-	20	24505900	0+2-	INS	-235	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24507963	3+1-	20	24508104	0+2-	INS	-140	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24519316	3+2-	20	24519301	3+2-	INS	-397	21	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	24521222	2+2-	20	24521213	2+2-	INS	-235	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	24548130	2+4-	20	24548160	2+4-	INS	-109	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24549698	3+3-	20	24549724	3+3-	INS	-179	29	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24577669	3+3-	20	24577656	3+3-	INS	-286	36	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24589998	3+0-	20	24590150	1+9-	INS	-149	29	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	24590137	4+0-	20	24590150	0+5-	INS	-185	29	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	24592636	2+0-	20	24592715	0+2-	INS	-245	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24610768	5+0-	20	24611194	1+3-	DEL	83	45	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24610768	3+0-	20	24610774	0+5-	DEL	93	49	3	COLO-829BL-IL|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	24612812	2+0-	20	24612911	0+2-	INS	-221	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24638223	3+3-	20	24638241	3+3-	INS	-373	30	3	COLO-829_v2_74|3	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24667617	2+3-	20	24667619	2+3-	INS	-118	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24679486	4+2-	20	24679521	4+2-	INS	-393	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24693483	3+0-	20	24693527	0+3-	INS	-277	37	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	24693997	2+3-	20	24693993	2+3-	INS	-394	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24700840	5+6-	20	24700821	5+6-	INS	-102	81	5	COLO-829BL-IL|1:COLO-829-IL|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	24721299	2+2-	20	24721318	2+2-	INS	-250	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24722367	6+5-	20	24722377	6+5-	INS	-91	71	5	COLO-829BL-IL|2:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24729693	4+1-	20	24729774	0+3-	INS	-202	42	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	24735891	2+6-	20	24736031	2+6-	INS	-273	11	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24748960	2+2-	20	24748968	2+2-	INS	-250	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24754023	2+1-	20	24754149	0+2-	INS	-195	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24764828	2+2-	20	24764876	2+2-	INS	-88	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24783659	2+2-	20	24783651	2+2-	INS	-110	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24789238	2+3-	20	24789294	2+3-	INS	-94	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24792326	2+2-	20	24792272	2+2-	INS	-265	32	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24804423	2+2-	20	24804404	2+2-	INS	-239	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24819085	4+1-	20	24819139	1+4-	INS	-202	54	5	COLO-829_v2_74|3:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	24821524	2+0-	20	24821928	0+3-	DEL	78	56	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	24821684	6+0-	20	24821696	1+5-	DEL	90	86	5	COLO-829BL-IL|3:COLO-829-IL|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	24842204	3+1-	20	24842286	0+3-	DEL	90	40	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24851715	14+1-	20	24852434	1+11-	DEL	725	99	11	COLO-829BL-IL|1:COLO-829-IL|10	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	24863787	2+3-	20	24863800	2+3-	INS	-107	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24869052	2+1-	20	24869081	0+2-	INS	-276	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24873196	4+2-	20	24873236	4+2-	INS	-249	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	24892431	2+2-	20	24892452	2+2-	INS	-251	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	24905537	2+2-	20	24905535	2+2-	INS	-97	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24910914	6+0-	20	24910971	0+7-	DEL	97	87	5	COLO-829BL-IL|1:COLO-829-IL|4	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	24924092	3+0-	20	24924129	1+4-	INS	-220	43	4	COLO-829_v2_74|3:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	24934662	2+2-	20	24934619	2+2-	INS	-392	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24970148	2+0-	20	24970310	2+2-	INS	-119	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24970462	2+0-	20	24970478	0+2-	INS	-252	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24982600	2+0-	20	24982661	0+3-	INS	-226	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24983134	2+3-	20	24983105	2+3-	INS	-90	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	24989321	2+2-	20	24989299	2+2-	INS	-394	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	24995730	5+0-	20	24995726	6+14-	INS	-107	45	5	COLO-829_v2_74|1:COLO-829-IL|4	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	24995981	2+6-	20	24995964	0+4-	INS	-306	10	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25001714	2+4-	20	25001709	2+4-	INS	-107	27	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25022241	2+2-	20	25022214	2+2-	INS	-104	35	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25027903	2+3-	20	25027915	2+3-	INS	-123	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25035066	2+2-	20	25035035	2+2-	INS	-107	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25061304	2+2-	20	25061286	2+2-	INS	-368	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25072833	4+3-	20	25072862	4+3-	INS	-95	38	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25078458	2+0-	20	25078485	2+4-	INS	-214	31	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	25079816	3+2-	20	25079813	3+2-	INS	-107	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	25094053	2+0-	20	25094060	0+3-	INS	-300	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25099403	3+3-	20	25099425	3+3-	INS	-98	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25104655	3+0-	20	25104774	0+3-	INS	-203	36	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25109853	4+3-	20	25109855	4+3-	INS	-105	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25123001	2+1-	20	25123035	0+2-	INS	-298	21	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25130008	4+1-	20	25130082	0+3-	INS	-174	36	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25146402	82+81-	20	25146755	82+81-	INS	-184	99	46	COLO-829BL-IL|9:COLO-829_v2_74|15:COLO-829-IL|22	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	25158091	2+3-	20	25158063	2+3-	INS	-246	26	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25173989	3+1-	20	25174078	0+3-	INS	-202	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25197426	3+3-	20	25197447	3+3-	INS	-115	24	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	25222162	2+2-	20	25222166	2+2-	INS	-226	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25235364	2+2-	20	25235508	0+2-	INS	-153	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25248433	2+0-	20	25248542	0+2-	INS	-212	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25266445	3+0-	20	25266426	0+3-	INS	-213	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25267978	2+2-	20	25267955	2+2-	INS	-103	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	25315873	3+2-	20	25315893	3+2-	INS	-108	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25318246	3+3-	20	25318303	3+3-	INS	-275	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25321522	3+0-	20	25321613	6+2-	INS	-222	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25347089	2+2-	20	25347068	2+2-	INS	-103	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25356177	2+2-	20	25356235	0+2-	INS	-249	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25378052	2+5-	20	25378066	2+5-	INS	-124	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25396298	4+2-	20	25396362	0+2-	INS	-149	32	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25397143	0+7-	20	25397674	6+0-	ITX	363	99	6	COLO-829-IL|6	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	25397502	3+0-	20	25397975	0+2-	DEL	431	41	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25410333	2+0-	20	25410510	0+2-	INS	-150	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25416633	2+0-	20	25416642	0+2-	INS	-273	17	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25433584	2+2-	20	25433597	2+2-	INS	-88	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	25442965	2+2-	20	25442943	2+2-	INS	-372	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25446301	2+2-	20	25446296	2+2-	INS	-254	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	25452039	3+2-	20	25452034	3+2-	INS	-108	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25462622	2+3-	20	25462623	2+3-	INS	-386	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25475058	3+3-	20	25475106	3+3-	INS	-102	34	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25480410	3+1-	20	25480428	0+3-	INS	-254	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25493812	2+3-	20	25493799	2+3-	INS	-106	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25509398	2+4-	20	25509395	2+4-	INS	-378	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25521250	2+2-	20	25521224	2+2-	INS	-124	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25530398	17+16-	20	25530546	0+4-	INS	-104	99	14	COLO-829BL-IL|2:COLO-829_v2_74|2:COLO-829-IL|10	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	25530543	3+2-	20	25530546	0+2-	INS	-322	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25531082	8+0-	20	25531678	2+11-	DEL	347	99	8	COLO-829_v2_74|8	0.22	BreakDancerMax-0.0.1r81	|q10|o20
20	25535985	3+2-	20	25535995	3+2-	INS	-109	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25540747	2+2-	20	25540759	2+2-	INS	-222	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25550009	2+0-	20	25550062	1+2-	INS	-270	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25554162	3+1-	20	25554228	3+6-	INS	-124	39	5	COLO-829BL-IL|2:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25555833	2+2-	20	25555789	2+2-	INS	-270	28	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25571082	2+3-	20	25571078	2+3-	INS	-102	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25595683	2+3-	20	25595676	2+3-	INS	-115	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25596691	2+1-	20	25596852	0+3-	INS	-142	21	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	25628454	2+2-	20	25628476	2+2-	INS	-103	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	25634961	2+4-	20	25634998	2+4-	INS	-95	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25646738	2+1-	20	25646825	2+3-	INS	-247	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25660600	2+2-	20	25660611	2+2-	INS	-104	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25666222	4+2-	20	25666211	4+2-	INS	-94	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25685935	35+14-	20	25686164	35+14-	INS	-95	25	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25689804	41+19-	20	25690038	41+19-	INS	-127	16	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25722291	12+1-	20	25784259	8+22-	DEL	61951	99	12	COLO-829BL-IL|4:COLO-829-IL|8	0.57	BreakDancerMax-0.0.1r81	|q10|o20
20	25778479	2+3-	20	25778535	2+3-	INS	-94	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	25785000	3+4-	20	25792225	12+1-	ITX	7103	51	3	COLO-829BL-IL|1:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25785899	2+13-	20	25793070	14+26-	ITX	7103	99	7	COLO-829BL-IL|3:COLO-829-IL|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25786172	5+2-	20	25796077	1+13-	DEL	9924	55	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25788602	1+2-	20	25796605	4+0-	ITX	7810	43	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25789897	4+7-	20	25791329	9+0-	ITX	1254	99	7	COLO-829BL-IL|1:COLO-829-IL|6	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	25789897	4+0-	20	25791573	0+3-	DEL	1654	64	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25815771	25+5-	20	25815820	25+5-	INS	-108	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25825187	59+1-	20	25825276	3+9-	INS	-199	10	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25832747	133+39-	20	25832921	133+39-	INS	-94	99	20	COLO-829BL-IL|5:COLO-829-IL|15	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	25833388	14+55-	20	25833497	14+55-	INS	-95	29	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25860458	2+2-	20	25860454	2+2-	INS	-114	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25886352	2+8-	20	25886340	2+8-	INS	-97	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25888080	5+43-	20	25888309	5+9-	INS	-110	13	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25897250	2+2-	20	25897258	2+2-	INS	-89	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25897781	2+2-	20	25897752	2+2-	ITX	-125	51	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25681477	45+34-	20	26032026	10+1-	INV	350553	99	7	COLO-829-IL|7	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25681477	37+33-	20	26032264	2+48-	INV	350797	81	3	COLO-829BL-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25681691	3+42-	20	26031666	3+24-	INV	349894	77	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25683621	1+12-	20	26030003	1+21-	INV	346345	99	9	COLO-829BL-IL|4:COLO-829-IL|5	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	25683922	38+10-	20	26029382	33+5-	INV	345436	99	25	COLO-829BL-IL|11:COLO-829-IL|14	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	25683922	12+9-	20	26029698	2+10-	INV	345747	99	7	COLO-829BL-IL|3:COLO-829-IL|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25685441	6+7-	20	26028182	4+170-	INV	342617	50	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25685872	2+8-	20	26027488	2+3-	INV	341495	62	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25686234	32+11-	20	26027156	28+19-	INV	340882	99	5	COLO-829_v2_74|4:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25686234	27+11-	20	26027648	32+26-	INV	341584	99	8	COLO-829BL-IL|5:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25686759	3+12-	20	26026660	48+43-	INV	339884	46	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25686970	18+22-	20	26026660	45+42-	INV	339599	99	13	COLO-829BL-IL|6:COLO-829-IL|7	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	25687768	0+2-	20	26025850	58+12-	INV	337983	55	2	COLO-829BL-IL|1:COLO-829-IL|1	0.20	BreakDancerMax-0.0.1r81	|q10|o20
20	25688354	19+20-	20	26025110	14+8-	INV	336745	99	7	COLO-829BL-IL|2:COLO-829-IL|5	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25688354	12+20-	20	26025339	0+3-	INV	336899	44	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25689098	2+0-	20	26024265	2+1-	INV	335053	59	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25691706	5+36-	20	26022177	8+47-	INV	330375	99	36	COLO-829BL-IL|14:COLO-829-IL|22	0.33	BreakDancerMax-0.0.1r81	|q10|o20
20	25691706	5+0-	20	26021948	6+0-	INV	330122	99	5	COLO-829BL-IL|1:COLO-829-IL|4	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	25692983	3+1-	20	26020684	4+3-	INV	327604	53	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25702325	23+35-	20	26011585	1+18-	INV	309177	99	18	COLO-829BL-IL|5:COLO-829-IL|13	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	25702776	16+2-	20	26010927	5+0-	INV	308091	86	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25703570	13+12-	20	26010048	3+0-	INV	306363	74	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25703570	10+12-	20	26010368	0+2-	INV	306744	59	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25703570	10+10-	20	26010131	2+1-	INV	306540	56	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25704243	58+27-	20	26009714	4+40-	INV	305467	99	19	COLO-829BL-IL|9:COLO-829-IL|10	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	25704243	58+8-	20	26009004	51+37-	INV	304757	99	30	COLO-829BL-IL|7:COLO-829-IL|23	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	25704243	28+8-	20	26009292	0+4-	INV	304948	72	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25704473	6+53-	20	26009004	21+37-	INV	304628	99	14	COLO-829BL-IL|3:COLO-829-IL|11	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	25937814	2+0-	20	25937989	0+5-	INS	-155	14	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	26023228	6+0-	20	26023628	0+2-	DEL	77	57	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26031148	15+10-	20	26031162	15+10-	INS	-102	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26075547	3+8-	20	26075599	3+8-	INS	-97	36	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	26077237	35+30-	20	26077292	35+30-	INS	-94	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26086439	5+9-	20	26086455	5+9-	INS	-115	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26092521	6+2-	20	26092533	6+2-	INS	-99	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26095212	99+66-	20	26095416	99+66-	INS	-92	23	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26097057	32+28-	20	26097305	16+47-	DEL	301	99	14	COLO-829BL-IL|7:COLO-829_v2_74|1:COLO-829-IL|6	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	26104305	2+2-	20	26104252	2+2-	INS	-113	37	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26105043	2+2-	20	26105037	2+2-	INS	-246	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26105967	3+3-	20	26105946	3+3-	INS	-283	35	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26136881	5+3-	20	26136893	5+3-	INS	-386	18	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26137034	9+10-	20	26137126	9+10-	INS	-96	99	9	COLO-829BL-IL|3:COLO-829-IL|6	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26138010	17+15-	20	26138238	17+15-	INS	-198	42	6	COLO-829BL-IL|2:COLO-829_v2_74|2:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26143128	2+2-	20	26143110	2+2-	INS	-109	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26146389	2+0-	20	26146454	0+2-	INS	-270	27	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	26148829	9+4-	20	26148822	9+4-	INS	-115	45	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26149671	43+12-	20	26149669	3+97-	INS	-290	8	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26151960	2+0-	20	26151944	142+23-	INS	-177	24	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	26152349	52+91-	20	26152482	52+91-	INS	-108	18	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26153888	52+27-	20	26154092	52+27-	INS	-252	11	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26154221	15+3-	20	26154203	15+3-	INS	-93	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26156567	7+53-	20	26156615	7+53-	INS	-108	26	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26157524	18+7-	20	26157607	18+7-	INS	-97	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26158486	5+3-	20	26158497	5+3-	ITX	-124	45	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26158736	12+0-	20	26158989	164+8-	INS	-91	45	4	COLO-829BL-IL|3:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26158915	45+12-	20	26158989	158+4-	INV	1	99	45	COLO-829BL-IL|17:COLO-829-IL|28	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	25807028	23+8-	20	26200385	5+10-	INV	393325	99	6	COLO-829BL-IL|2:COLO-829-IL|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25807163	24+8-	20	26199924	79+33-	INV	392701	99	20	COLO-829BL-IL|8:COLO-829-IL|12	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	25807163	4+8-	20	26200146	3+26-	INV	392956	99	7	COLO-829BL-IL|1:COLO-829-IL|6	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25807697	50+10-	20	26199609	16+10-	INV	391879	68	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25807697	50+7-	20	26199420	39+7-	INV	391725	99	26	COLO-829BL-IL|7:COLO-829-IL|19	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	25808397	2+3-	20	26198892	11+9-	INV	390472	48	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	25808510	34+2-	20	26198892	11+7-	INV	390280	48	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25808510	34+0-	20	26198477	18+30-	INV	389994	99	7	COLO-829BL-IL|3:COLO-829-IL|4	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	25808846	44+34-	20	26198477	10+29-	INV	389579	99	19	COLO-829BL-IL|8:COLO-829-IL|11	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	25809924	5+1-	20	26197102	11+7-	INV	387089	47	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25810501	7+38-	20	26196849	34+29-	INV	386265	99	27	COLO-829BL-IL|11:COLO-829-IL|16	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	25810971	14+9-	20	26196064	10+17-	INV	385141	99	7	COLO-829-IL|7	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	25810971	7+9-	20	26196300	2+14-	INV	385246	99	7	COLO-829BL-IL|4:COLO-829-IL|3	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	25813421	2+0-	20	26193337	3+0-	INV	379588	70	2	COLO-829_v2_74|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	25813562	6+0-	20	26193438	7+2-	INV	379719	99	6	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|3	0.21	BreakDancerMax-0.0.1r81	|q10|o20
20	25814186	1+2-	20	26193438	1+2-	INV	378900	66	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25815890	23+3-	20	26191425	14+2-	INV	375539	47	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25818260	9+6-	20	26189063	7+17-	INV	370833	92	4	COLO-829BL-IL|2:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25818260	9+2-	20	26188847	4+2-	INV	370584	42	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25818837	18+10-	20	26188491	0+7-	INV	369614	99	7	COLO-829BL-IL|4:COLO-829-IL|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	25819074	14+6-	20	26187998	6+1-	INV	368822	99	6	COLO-829BL-IL|2:COLO-829-IL|4	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	25820267	3+17-	20	26186904	3+0-	INV	366602	84	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	25821011	2+5-	20	26186358	2+4-	INV	365264	52	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	26162342	6+0-	20	26168365	4+39-	INS	-101	19	2	COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	26181376	11+3-	20	26181479	2+28-	DEL	95	99	11	COLO-829BL-IL|7:COLO-829-IL|4	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	26187063	2+2-	20	26187025	2+2-	INS	-108	33	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	25803321	8+5-	20	26203624	7+6-	INV	400240	99	6	COLO-829BL-IL|3:COLO-829-IL|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	25804441	9+8-	20	26202591	10+18-	INV	398179	99	6	COLO-829BL-IL|2:COLO-829-IL|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25805083	9+11-	20	26201834	34+19-	INV	396860	99	9	COLO-829BL-IL|4:COLO-829-IL|5	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	25805083	0+11-	20	26202256	8+27-	INV	397072	99	9	COLO-829BL-IL|2:COLO-829-IL|7	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	25805546	15+33-	20	26201834	25+19-	INV	396229	87	4	COLO-829BL-IL|1:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	25805764	13+9-	20	26201291	59+32-	INV	395508	99	13	COLO-829BL-IL|3:COLO-829-IL|10	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	25805764	0+9-	20	26201594	0+10-	INV	395780	99	9	COLO-829BL-IL|3:COLO-829-IL|6	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	25806681	3+34-	20	26200623	20+59-	INV	393884	99	33	COLO-829BL-IL|14:COLO-829-IL|19	0.42	BreakDancerMax-0.0.1r81	|q10|o20
20	26185682	21+23-	20	26204340	1+2-	INV	18551	43	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26185682	20+20-	20	26204005	18+19-	INV	18281	99	17	COLO-829BL-IL|6:COLO-829-IL|11	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	26203157	4+2-	20	26203111	4+2-	INS	-121	36	2	COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	26207055	112+95-	20	26207139	0+5-	DEL	91	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26207586	5+4-	20	26207578	2+3-	INS	-298	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26209421	6+4-	20	26209427	6+4-	INS	-245	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26213026	35+21-	20	26216063	27+24-	DEL	3014	99	11	COLO-829BL-IL|7:COLO-829-IL|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	26216165	27+13-	20	26223162	41+37-	ITX	6971	99	7	COLO-829BL-IL|4:COLO-829-IL|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	26222016	36+21-	20	26223162	34+37-	ITX	842	62	4	COLO-829BL-IL|3:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26216300	7+5-	20	26223455	2+1-	ITX	6961	42	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26220407	57+14-	20	26220546	11+9-	DEL	92	86	4	COLO-829BL-IL|2:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26221124	2+2-	20	26221077	2+2-	INS	-110	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26222442	3+2-	20	26222442	3+2-	INS	-100	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26213026	24+21-	20	26228746	7+24-	DEL	15857	46	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26213026	21+21-	20	26234778	2+6-	DEL	21734	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26213026	19+21-	20	26227865	2+3-	DEL	14801	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26222016	35+17-	20	26228746	7+21-	DEL	6926	56	4	COLO-829BL-IL|2:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26234763	15+6-	20	26234778	2+4-	DEL	89	34	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26216300	7+3-	20	26250275	9+28-	DEL	33933	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26223417	31+37-	20	26250275	9+26-	DEL	26914	99	12	COLO-829BL-IL|6:COLO-829-IL|6	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	26235284	76+33-	20	26235304	14+49-	DEL	88	43	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26236941	4+1-	20	26237002	47+27-	DEL	90	47	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26237570	13+11-	20	26237748	13+11-	INS	-196	20	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26238514	6+2-	20	26238580	1+4-	DEL	91	56	3	COLO-829BL-IL|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	26245212	22+20-	20	26245237	1+2-	INS	-292	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26246991	4+2-	20	26246986	10+13-	INS	-160	21	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26247155	9+10-	20	26248537	18+56-	DEL	1204	64	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26247458	53+36-	20	26248537	18+53-	DEL	1200	99	39	COLO-829BL-IL|13:COLO-829-IL|26	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	26249703	12+14-	20	26253640	391+278-	INS	-109	44	4	COLO-829BL-IL|1:COLO-829-IL|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	26253795	385+274-	20	26253852	19+18-	DEL	89	99	6	COLO-829BL-IL|3:COLO-829-IL|3	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26250981	6+2-	20	26250999	6+2-	INS	-110	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26251219	4+0-	20	26251213	55+59-	ITX	-147	36	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26256261	13+6-	20	26256321	13+6-	INS	-195	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26210853	13+4-	20	26263379	12+86-	DEL	52506	42	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26221388	12+15-	20	26263379	12+84-	DEL	41976	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26263509	12+82-	20	26263543	32+18-	DEL	90	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26261120	490+169-	20	26263379	10+82-	DEL	2286	99	8	COLO-829BL-IL|2:COLO-829-IL|6	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26253795	379+274-	20	26263379	10+74-	DEL	9591	99	10	COLO-829BL-IL|5:COLO-829-IL|5	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26261572	58+42-	20	26263379	10+64-	DEL	1917	60	4	COLO-829BL-IL|2:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26249703	12+12-	20	26263543	31+15-	DEL	13877	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	26260002	22+82-	20	26260842	482+169-	DEL	1063	53	4	COLO-829BL-IL|1:COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26261120	482+165-	20	26262210	19+54-	ITX	975	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26252375	69+32-	20	26260842	482+163-	DEL	8713	40	3	COLO-829BL-IL|1:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26261120	482+160-	20	26261252	54+42-	DEL	89	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26253795	369+274-	20	26262210	17+54-	DEL	8409	35	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26253795	367+274-	20	26259671	17+81-	DEL	5996	99	12	COLO-829BL-IL|5:COLO-829-IL|7	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26260002	17+69-	20	26261974	24+9-	ITX	1298	41	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26252375	65+31-	20	26263063	16+25-	DEL	10775	99	7	COLO-829BL-IL|5:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26245212	20+20-	20	26265972	83+122-	DEL	20859	82	5	COLO-829BL-IL|1:COLO-829-IL|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	26266174	83+117-	20	26267368	32+50-	ITX	1142	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26266174	83+115-	20	26266365	93+253-	DEL	85	99	8	COLO-829BL-IL|2:COLO-829_v2_74|3:COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26265954	12+10-	20	26265972	80+114-	DEL	93	59	4	COLO-829BL-IL|1:COLO-829-IL|3	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26266366	105+125-	20	26266365	84+242-	DEL	97	99	26	COLO-829BL-IL|14:COLO-829-IL|12	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26265480	39+46-	20	26266365	84+216-	ITX	940	38	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	26266786	81+216-	20	26266768	7+9-	DEL	93	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	26265075	11+10-	20	26265197	38+42-	DEL	159	99	7	COLO-829BL-IL|1:COLO-829-IL|6	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	28034669	15+7-	20	28034766	15+7-	INS	-199	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28047791	7+9-	20	28047864	7+9-	INS	-94	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28048396	4+5-	20	28048442	9+14-	DEL	148	96	6	COLO-829BL-IL|1:COLO-829-IL|5	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	28054182	13+5-	20	28054205	13+5-	INS	-221	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28054708	65+95-	20	28055961	6+10-	DEL	1308	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28055281	2+2-	20	28055264	2+2-	INS	-99	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28061931	6+4-	20	28061908	6+4-	INS	-102	64	4	COLO-829BL-IL|1:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	28069549	5+15-	20	28069582	5+15-	INS	-93	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28083852	10+2-	20	28083908	10+2-	INS	-114	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28086059	34+1-	20	28087210	5+28-	DEL	1150	99	23	COLO-829BL-IL|6:COLO-829-IL|17	0.21	BreakDancerMax-0.0.1r81	|q10|o20
20	28091892	2+3-	20	28091939	2+3-	INS	-106	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28099587	27+4-	20	28099640	27+4-	INS	-93	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28111198	20+8-	20	28111288	20+8-	INS	-245	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28131579	5+1-	20	28131583	0+3-	INS	-93	51	3	COLO-829BL-IL|1:COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	28155101	9+17-	20	28155205	9+17-	INS	-107	18	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28181031	2+2-	20	28181037	2+2-	INS	-103	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28190139	11+2-	20	28190136	11+2-	INS	-230	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	28195773	56+34-	20	28195962	56+34-	ITX	-129	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28196681	458+69-	20	28197332	458+69-	INS	-141	21	5	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28199206	20+13-	20	28199202	20+13-	INS	-109	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28200289	197+13-	20	28200440	197+13-	INS	-105	16	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28201703	189+243-	20	28202001	189+243-	INS	-102	13	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28203851	238+33-	20	28203967	238+33-	INS	-105	22	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28204578	3+47-	20	28204638	0+11-	INS	-190	14	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28205445	6+3-	20	28205508	6+3-	INS	-102	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28206055	16+40-	20	28206247	16+40-	INS	-126	16	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28207096	136+176-	20	28207397	136+176-	INS	-103	12	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28207920	8+33-	20	28208006	8+33-	INS	-108	30	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28208829	18+32-	20	28209678	7+23-	DEL	897	99	12	COLO-829BL-IL|3:COLO-829-IL|9	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	28209189	241+119-	20	28209623	241+119-	INS	-108	11	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28213322	3+10-	20	28213337	8+5-	INS	-240	33	4	COLO-829_v2_74|3:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28214448	52+51-	20	28214718	52+51-	INS	-107	14	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28221074	11+244-	20	28221129	11+244-	INS	-230	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28221403	50+65-	20	28221813	50+65-	INS	-110	18	4	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28227059	55+33-	20	28227180	55+33-	INS	-99	22	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28227671	35+7-	20	28227701	35+7-	INS	-104	38	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	28229839	26+63-	20	28229889	26+63-	INS	-118	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28230042	94+6-	20	28230168	94+6-	INS	-116	18	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28230864	43+78-	20	28231023	43+78-	ITX	-130	30	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28231460	20+9-	20	28231439	20+9-	INS	-94	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28232599	53+112-	20	28232997	53+112-	INS	-107	26	4	COLO-829BL-IL|2:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28234680	188+73-	20	28234791	188+73-	INS	-178	23	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28234973	29+172-	20	28235130	29+172-	INS	-95	28	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28239389	306+354-	20	28239877	306+354-	INS	-113	9	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28240030	3+6-	20	28240040	3+6-	INS	-102	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28240366	7+19-	20	28240407	7+19-	INS	-94	36	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28242759	249+222-	20	28242753	110+16-	INS	-187	27	5	COLO-829_v2_74|4:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28243007	171+81-	20	28243133	171+81-	INS	-95	22	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28243326	304+243-	20	28243660	304+243-	INS	-99	99	49	COLO-829BL-IL|17:COLO-829-IL|32	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	28243853	22+84-	20	28243869	22+84-	INS	-246	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28244745	48+558-	20	28244826	48+558-	INS	-99	33	3	COLO-829BL-IL|2:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28245559	27+55-	20	28245959	27+55-	INS	-92	11	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28246268	9+179-	20	28246479	9+179-	INS	-104	25	3	COLO-829BL-IL|2:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28247503	215+232-	20	28247689	215+232-	INS	-123	24	3	COLO-829BL-IL|1:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28248243	973+726-	20	28249058	973+726-	INS	-121	40	9	COLO-829BL-IL|3:COLO-829_v2_74|2:COLO-829-IL|4	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28249464	186+455-	20	28250381	186+455-	INS	-125	97	16	COLO-829BL-IL|2:COLO-829_v2_74|3:COLO-829-IL|11	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28250690	846+675-	20	28252461	846+675-	INS	-148	99	37	COLO-829BL-IL|9:COLO-829_v2_74|11:COLO-829-IL|17	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28252531	808+637-	20	28255183	113+276-	DEL	971	99	20	COLO-829BL-IL|6:COLO-829_v2_74|7:COLO-829-IL|7	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28252531	801+637-	20	28255064	41+88-	DEL	2599	99	86	COLO-829BL-IL|37:COLO-829_v2_74|2:COLO-829-IL|47	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28252961	2+2-	20	28252942	2+2-	INS	-100	29	2	COLO-829-IL|2	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	28259691	8+28-	20	28259840	8+28-	INS	-104	16	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28259910	6+26-	20	28259893	43+52-	DEL	90	99	22	COLO-829BL-IL|8:COLO-829_v2_74|1:COLO-829-IL|13	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28260476	11+16-	20	28260472	14+10-	INS	-154	15	4	COLO-829_v2_74|1:COLO-829-IL|3	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28260768	10+3-	20	28260754	92+19-	INS	-157	26	6	COLO-829BL-IL|2:COLO-829_v2_74|3:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28261160	89+13-	20	28261146	13+51-	DEL	95	99	47	COLO-829BL-IL|14:COLO-829_v2_74|6:COLO-829-IL|27	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	28261160	41+13-	20	28261620	12+69-	DEL	211	99	24	COLO-829_v2_74|24	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28261579	12+2-	20	28261620	7+40-	DEL	95	99	12	COLO-829BL-IL|4:COLO-829_v2_74|4:COLO-829-IL|4	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	28262622	9+6-	20	28262670	9+6-	INS	-113	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28263313	105+225-	20	28264009	105+225-	INS	-163	43	10	COLO-829BL-IL|3:COLO-829_v2_74|6:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28264227	168+119-	20	28265145	168+119-	INS	-156	71	14	COLO-829BL-IL|6:COLO-829_v2_74|4:COLO-829-IL|4	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28265505	216+15-	20	28265881	216+15-	INS	-123	74	10	COLO-829BL-IL|4:COLO-829_v2_74|2:COLO-829-IL|4	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28266051	13+108-	20	28266251	13+108-	INS	-146	42	5	COLO-829BL-IL|3:COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28266480	58+13-	20	28266544	58+13-	INS	-255	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	28266694	746+99-	20	28267531	746+99-	INS	-214	19	7	COLO-829BL-IL|1:COLO-829_v2_74|4:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	29267646	38+36-	20	29267622	38+36-	INS	-98	99	15	COLO-829BL-IL|4:COLO-829-IL|11	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	29268290	20+6-	20	29268646	4+2-	DEL	78	40	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29268290	18+6-	20	29268377	7+21-	INS	-139	15	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29268789	4+0-	20	29269013	5+11-	DEL	76	40	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29268996	24+18-	20	29269013	5+9-	DEL	89	80	5	COLO-829BL-IL|4:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29269322	5+4-	20	29269352	2+4-	INS	-273	9	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29269843	10+2-	20	29270092	42+68-	DEL	84	99	12	COLO-829BL-IL|2:COLO-829_v2_74|6:COLO-829-IL|4	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	29270447	36+56-	20	29270645	1+4-	DEL	77	84	4	COLO-829_v2_74|4	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29273620	5+3-	20	29273630	3+6-	INS	-187	11	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29274378	27+23-	20	29274639	9+8-	INS	-165	21	5	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29275073	9+6-	20	29275143	0+3-	INS	-114	21	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29275681	256+189-	20	29275914	459+444-	DEL	91	99	283	COLO-829BL-IL|154:COLO-829_v2_74|1:COLO-829-IL|128	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	29275681	242+177-	20	29279248	156+115-	DEL	3252	63	3	COLO-829_v2_74|3	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	29275681	239+177-	20	29275687	18+22-	DEL	89	94	6	COLO-829BL-IL|4:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	29276711	152+135-	20	29276730	35+26-	INS	-191	3	3	COLO-829_v2_74|2:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	29275913	18+15-	20	29275914	150+135-	DEL	89	99	11	COLO-829BL-IL|2:COLO-829-IL|9	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	29278877	11+2-	20	29279248	156+112-	DEL	78	99	6	COLO-829_v2_74|6	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	29279378	156+106-	20	29279761	5+25-	DEL	77	99	12	COLO-829_v2_74|12	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	29277142	32+21-	20	29277464	15+30-	DEL	78	99	12	COLO-829_v2_74|12	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29279466	14+9-	20	29279761	4+12-	DEL	77	99	8	COLO-829_v2_74|8	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	29278988	20+23-	20	29279362	6+9-	DEL	77	79	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29275681	232+177-	20	29292781	955+875-	DEL	238	99	233	COLO-829BL-IL|105:COLO-829_v2_74|11:COLO-829-IL|117	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	29293644	603+519-	20	29293651	44+69-	DEL	77	99	36	COLO-829_v2_74|36	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	29293644	567+519-	20	29293763	12+16-	DEL	78	99	6	COLO-829_v2_74|6	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	29293644	561+519-	20	29293968	22+22-	DEL	78	67	4	COLO-829_v2_74|4	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	29292169	20+19-	20	29292453	4+12-	DEL	79	38	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29286866	68+59-	20	29292453	4+10-	DEL	988	99	12	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|9	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29294260	20+16-	20	29294519	5+11-	DEL	77	99	5	COLO-829_v2_74|5	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29294260	15+16-	20	29294677	21+21-	DEL	78	36	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	29291956	11+1-	20	29291937	17+18-	DEL	88	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29291606	3+5-	20	29291937	17+15-	DEL	78	41	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29286177	6+4-	20	29286383	47+40-	DEL	77	35	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29286866	47+38-	20	29286856	0+11-	DEL	90	99	11	COLO-829BL-IL|6:COLO-829-IL|5	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29294371	11+5-	20	29294677	21+19-	DEL	77	90	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29294982	21+15-	20	29295208	8+4-	DEL	77	40	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29291150	52+42-	20	29291448	1+5-	DEL	77	99	5	COLO-829_v2_74|5	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29285595	37+21-	20	29285959	4+4-	DEL	83	56	4	COLO-829_v2_74|2:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29295351	8+2-	20	29295659	35+49-	DEL	78	99	6	COLO-829_v2_74|6	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	29290582	8+1-	20	29290790	46+41-	DEL	78	99	6	COLO-829_v2_74|6	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29285595	31+17-	20	29285577	16+49-	DEL	82	55	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29295571	8+3-	20	29295659	35+43-	DEL	91	57	4	COLO-829BL-IL|1:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29285777	16+44-	20	29285785	2+6-	INS	-267	10	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29285777	12+44-	20	29286168	0+2-	DEL	78	46	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29280889	14+19-	20	29281156	9+5-	DEL	77	40	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29281433	9+3-	20	29281425	125+92-	INS	-176	9	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29281791	123+86-	20	29281959	0+6-	DEL	77	99	6	COLO-829_v2_74|6	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29281791	117+86-	20	29282025	46+33-	DEL	78	99	7	COLO-829_v2_74|7	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29281036	38+10-	20	29281425	110+86-	DEL	78	99	27	COLO-829_v2_74|27	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	29282332	46+26-	20	29282577	14+15-	DEL	77	99	8	COLO-829_v2_74|8	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29283319	4+3-	20	29283303	6+7-	INS	-262	9	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29283518	6+5-	20	29283874	1+6-	DEL	78	45	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29283693	6+0-	20	29284077	7+9-	DEL	77	99	6	COLO-829_v2_74|6	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	29284250	7+3-	20	29284619	15+7-	DEL	78	41	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29288568	13+3-	20	29288956	3+6-	DEL	77	99	4	COLO-829_v2_74|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	29289097	3+2-	20	29289390	7+13-	DEL	78	46	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29289545	7+11-	20	29289953	4+5-	DEL	77	41	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29296032	16+15-	20	29296162	16+15-	INS	-95	95	8	COLO-829BL-IL|4:COLO-829-IL|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29310545	2+2-	20	29310530	2+2-	INS	-88	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29323251	2+2-	20	29323229	2+2-	INS	-120	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29353880	3+2-	20	29353933	3+2-	INS	-107	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29376815	2+2-	20	29376785	2+2-	INS	-380	24	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	29394102	4+3-	20	29394117	4+3-	INS	-109	41	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29404342	2+2-	20	29404355	2+2-	INS	-110	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	29405003	2+2-	20	29404959	2+2-	INS	-108	35	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29418954	2+0-	20	29419087	0+2-	INS	-174	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29424296	2+2-	20	29424249	2+2-	INS	-115	36	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29439173	2+2-	20	29439153	2+2-	INS	-90	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29449647	3+2-	20	29449626	3+2-	INS	-118	30	2	COLO-829-IL|2	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	29457801	4+4-	20	29457872	4+4-	INS	-216	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29459696	2+2-	20	29459664	2+2-	INS	-395	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29465146	3+1-	20	29465243	0+2-	INS	-224	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29466079	2+2-	20	29466068	2+2-	INS	-235	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29469066	2+2-	20	29469017	2+2-	INS	-110	37	2	COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	29471701	2+2-	20	29471649	2+2-	INS	-401	31	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29497730	2+2-	20	29497697	2+2-	INS	-95	36	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29504571	3+2-	20	29504549	3+2-	INS	-246	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29580585	2+0-	20	29580791	1+4-	INS	-106	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29586615	2+4-	20	29586652	2+4-	INS	-219	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29604310	2+2-	20	29604276	2+2-	INS	-384	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29627358	2+2-	20	29627312	2+2-	INS	-109	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	29643107	3+3-	20	29643181	3+3-	INS	-209	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29657894	2+1-	20	29657956	1+3-	INS	-210	40	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	29686036	2+3-	20	29686062	2+3-	INS	-90	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29697479	2+2-	20	29697523	2+2-	INS	-98	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29733284	2+2-	20	29733320	2+2-	INS	-230	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29737004	5+4-	20	29737009	5+4-	INS	-228	43	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	29740806	2+2-	20	29740822	2+2-	INS	-215	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29759420	2+3-	20	29759407	2+3-	INS	-118	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29762708	3+1-	20	29762796	1+3-	INS	-215	23	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29768929	2+2-	20	29768911	2+2-	INS	-375	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29771002	4+2-	20	29771020	4+2-	INS	-248	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29771090	2+0-	20	29771174	1+3-	INS	-274	21	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29772685	2+2-	20	29772645	2+2-	INS	-101	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29818816	2+3-	20	29818885	2+3-	INS	-102	21	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29857054	3+3-	20	29857091	3+3-	INS	-207	28	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29857761	2+2-	20	29857737	2+2-	INS	-103	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	29873823	2+0-	20	29873939	1+3-	INS	-173	30	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	29893843	2+2-	20	29893831	2+2-	INS	-232	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	29920608	4+3-	20	29920675	4+3-	INS	-197	30	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29939714	3+3-	20	29939760	3+3-	INS	-207	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	29941475	5+11-	20	29941459	5+11-	INS	-106	79	5	COLO-829BL-IL|2:COLO-829-IL|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	29946681	2+1-	20	29946855	0+2-	INS	-146	19	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	29986931	3+4-	20	29987019	3+4-	INS	-192	25	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30009585	3+2-	20	30009567	3+2-	ITX	-126	42	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30016371	3+3-	20	30016365	3+3-	INS	-387	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30016838	3+2-	20	30016861	3+2-	INS	-242	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30022828	2+0-	20	30023043	1+2-	INS	-123	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30024442	3+4-	20	30024477	3+4-	INS	-90	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30025937	2+0-	20	30025937	0+4-	INS	-288	14	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30032116	2+0-	20	30032189	1+2-	INS	-234	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30043105	3+3-	20	30043178	3+3-	INS	-93	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30053112	2+2-	20	30053089	2+2-	INS	-373	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30074913	2+2-	20	30074917	2+2-	INS	-87	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30077711	2+4-	20	30077751	2+4-	INS	-87	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	30091705	2+2-	20	30091692	2+2-	INS	-244	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	30096954	2+2-	20	30096978	2+2-	INS	-239	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30106688	4+4-	20	30106809	4+4-	INS	-257	28	4	COLO-829_v2_74|3:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30107167	2+2-	20	30107153	2+2-	INS	-109	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	30109192	2+2-	20	30109296	0+2-	INS	-189	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30114057	3+1-	20	30114050	1+4-	INS	-250	25	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	30130555	2+3-	20	30130619	2+3-	INS	-117	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30132654	2+0-	20	30132681	2+3-	INS	-209	30	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30134210	4+4-	20	30134236	4+4-	INS	-100	38	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30134746	2+3-	20	30134788	2+3-	INS	-211	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30145004	2+2-	20	30145015	2+2-	INS	-105	29	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	30149845	3+0-	20	30149963	1+2-	INS	-188	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30150199	2+4-	20	30150218	2+4-	INS	-109	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30150652	7+2-	20	30150703	7+2-	INS	-124	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30176536	2+2-	20	30176541	2+2-	INS	-104	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30177837	2+3-	20	30177792	2+3-	INS	-394	28	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30179068	2+1-	20	30179050	1+3-	INS	-323	23	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	30197188	3+4-	20	30197209	3+4-	INS	-301	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30200040	4+2-	20	30200041	4+2-	INS	-378	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30210052	3+4-	20	30210129	3+4-	INS	-95	24	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30238300	2+2-	20	30238246	2+2-	INS	-117	37	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30239441	2+3-	20	30239461	2+3-	INS	-376	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30240987	4+1-	20	30241185	0+3-	INS	-143	37	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30247000	2+2-	20	30247019	2+2-	INS	-331	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30261709	2+2-	20	30261715	2+2-	INS	-96	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30278411	2+2-	20	30278421	2+2-	INS	-216	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30288962	2+3-	20	30288975	2+3-	INS	-98	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30296697	2+2-	20	30296706	2+2-	INS	-91	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30302592	2+5-	20	30302656	2+5-	INS	-234	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30308741	4+5-	20	30308840	4+5-	INS	-175	37	4	COLO-829_v2_74|1:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30313959	3+1-	20	30314044	0+2-	INS	-161	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30314248	2+2-	20	30314239	2+2-	INS	-109	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30329886	4+1-	20	30329896	0+2-	INS	-271	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30361254	2+3-	20	30361292	2+3-	INS	-97	27	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30362563	4+1-	20	30363193	0+29-	DEL	314	99	4	COLO-829_v2_74|4	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	30362894	24+1-	20	30363193	0+25-	DEL	317	99	24	COLO-829BL-IL|5:COLO-829-IL|19	0.55	BreakDancerMax-0.0.1r81	|q10|o20
20	30370683	2+2-	20	30370660	2+2-	INS	-104	30	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	30382973	2+0-	20	30383088	2+2-	INS	-185	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30383187	2+0-	20	30383346	1+3-	INS	-141	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30401685	2+2-	20	30401650	2+2-	INS	-259	25	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30403823	2+1-	20	30403806	2+4-	INS	-251	23	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	30409088	2+2-	20	30409080	2+2-	INS	-257	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	30414930	2+3-	20	30414904	2+3-	INS	-244	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30434011	3+2-	20	30433971	3+2-	INS	-106	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30435542	2+0-	20	30435595	0+3-	INS	-281	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30455895	2+2-	20	30455913	2+2-	INS	-105	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30466416	2+2-	20	30466408	2+2-	INS	-112	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30470214	6+32-	20	30470294	6+32-	INS	-102	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30503499	2+2-	20	30503490	2+2-	INS	-100	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30530555	4+0-	20	30530580	0+3-	INS	-234	25	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	30540114	23+27-	20	30540458	23+27-	DEL	94	90	6	COLO-829BL-IL|1:COLO-829-IL|5	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30553672	2+2-	20	30553697	2+2-	INS	-104	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30562064	2+2-	20	30562079	2+2-	INS	-104	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30569760	2+2-	20	30569782	2+2-	INS	-113	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30597147	2+2-	20	30597092	2+2-	INS	-405	32	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30607238	2+2-	20	30607244	2+2-	INS	-93	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30609658	2+2-	20	30609670	2+2-	INS	-93	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30637828	2+2-	20	30637834	2+2-	INS	-101	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30680937	4+5-	20	30680986	4+5-	INS	-353	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30691920	2+0-	20	30693435	2+1-	INV	1408	57	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30708814	3+0-	20	30708904	2+3-	INS	-203	39	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	30709718	2+2-	20	30709700	2+2-	INS	-112	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30734181	3+1-	20	30734381	0+2-	INS	-110	37	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	30745516	2+2-	20	30745461	2+2-	INS	-113	39	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	30765214	2+3-	20	30765182	2+3-	INS	-116	36	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	30771269	2+2-	20	30771275	2+2-	INS	-96	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30774542	11+3-	20	30776412	0+15-	DEL	1913	99	11	COLO-829BL-IL|3:COLO-829-IL|8	0.35	BreakDancerMax-0.0.1r81	|q10|o20
20	30779869	2+2-	20	30779807	2+2-	INS	-122	44	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30786205	4+2-	20	30786267	4+2-	INS	-213	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30798622	2+2-	20	30798620	2+2-	INS	-111	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	30805052	2+2-	20	30805047	2+2-	INS	-241	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30807866	2+0-	20	30807877	0+2-	INS	-314	22	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	30828650	3+2-	20	30828670	3+2-	INS	-100	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30839681	2+2-	20	30839667	2+2-	INS	-228	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	30868870	4+3-	20	30868948	4+3-	INS	-105	20	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30877282	2+6-	20	30877288	2+6-	INS	-95	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30897707	2+2-	20	30897697	2+2-	INS	-108	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	30903248	2+2-	20	30903221	2+2-	INS	-98	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30909931	2+0-	20	30909916	0+2-	INS	-330	20	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	30914869	3+1-	20	30914885	0+2-	INS	-246	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	30916393	2+0-	20	30916591	0+2-	INS	-129	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30920833	3+3-	20	30920843	3+3-	INS	-99	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30953122	2+2-	20	30953109	2+2-	INS	-237	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30953905	2+0-	20	30954096	0+2-	INS	-143	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	30994762	2+2-	20	30994725	2+2-	INS	-399	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	30997656	2+0-	20	30997687	1+2-	INS	-240	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31044115	2+3-	20	31044086	2+3-	INS	-109	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31044663	2+2-	20	31044691	2+2-	INS	-97	24	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31046949	2+2-	20	31046945	2+2-	INS	-97	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31056280	2+2-	20	31056278	2+2-	INS	-237	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31075416	2+2-	20	31075375	2+2-	INS	-391	27	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31091335	2+2-	20	31091301	2+2-	INS	-103	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31092275	6+3-	20	31092385	6+3-	INS	-102	23	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31095133	2+2-	20	31095090	2+2-	INS	-393	27	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31098211	4+1-	20	31098286	0+2-	INS	-189	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31099364	2+2-	20	31099360	2+2-	INS	-114	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31101403	3+3-	20	31101430	3+3-	INS	-171	29	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31109129	3+7-	20	31109129	0+2-	INS	-89	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31115152	2+2-	20	31115148	2+2-	INS	-93	31	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31119088	2+2-	20	31119074	2+2-	INS	-235	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31137523	2+0-	20	31137592	0+3-	INS	-248	16	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	31139031	2+2-	20	31139038	2+2-	INS	-99	30	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31151639	2+1-	20	31151828	0+2-	INS	-117	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31161815	2+2-	20	31161758	2+2-	ITX	-130	54	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31163403	2+0-	20	31163504	0+2-	INS	-215	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31164662	2+2-	20	31164627	2+2-	INS	-108	36	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31183117	2+3-	20	31183088	2+3-	INS	-88	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31209023	2+0-	20	31209071	0+2-	INS	-265	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31242024	2+3-	20	31242034	2+3-	INS	-105	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31275645	2+3-	20	31275698	2+3-	INS	-88	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31297724	2+0-	20	31297719	0+3-	INS	-354	20	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	31300318	2+2-	20	31300257	2+2-	INS	-411	36	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31319669	3+2-	20	31319646	3+2-	INS	-100	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31334847	2+0-	20	31334975	0+2-	INS	-175	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31335994	2+0-	20	31336083	0+2-	INS	-226	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31355889	3+1-	20	31355875	0+2-	INS	-355	35	3	COLO-829_v2_74|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	31357412	2+0-	20	31357613	0+2-	INS	-131	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31377408	2+2-	20	31377401	2+2-	INS	-100	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31405159	2+2-	20	31405133	2+2-	INS	-95	35	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31406546	2+2-	20	31406565	2+2-	INS	-371	18	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	31411458	2+3-	20	31411507	2+3-	INS	-114	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31411900	2+2-	20	31411875	2+2-	INS	-86	34	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31414310	3+3-	20	31414310	3+3-	INS	-349	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31444931	2+2-	20	31444947	2+2-	INS	-101	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31455703	2+3-	20	31455741	2+3-	INS	-102	27	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31462436	2+2-	20	31462433	2+2-	INS	-221	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31465140	2+2-	20	31465130	2+2-	INS	-238	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31470787	2+4-	20	31470878	2+4-	INS	-223	15	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31496917	2+2-	20	31496878	2+2-	INS	-105	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31533954	3+1-	20	31533938	0+2-	INS	-99	38	3	COLO-829BL-IL|2:COLO-829-IL|1	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	31574507	3+1-	20	31574621	1+3-	INS	-164	41	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31580881	2+2-	20	31580880	2+2-	INS	-108	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31625169	2+2-	20	31625151	2+2-	INS	-89	33	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31645391	2+0-	20	31645381	2+2-	INS	-307	17	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	31645515	2+0-	20	31645538	1+2-	INS	-272	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31646147	2+0-	20	31646231	0+2-	INS	-242	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31647315	2+2-	20	31647280	2+2-	INS	-107	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31648094	2+2-	20	31648072	2+2-	INS	-372	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31686135	2+2-	20	31686188	2+2-	INS	-337	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31695663	2+3-	20	31695647	2+3-	INS	-93	33	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	31701918	4+4-	20	31702035	4+4-	INS	-189	23	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31728356	2+2-	20	31728316	2+2-	INS	-389	26	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31730910	2+2-	20	31730917	2+2-	INS	-96	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31733109	2+0-	20	31733297	1+2-	INS	-128	20	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	31756441	3+3-	20	31756479	3+3-	INS	-287	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	31763363	2+1-	20	31763448	0+3-	INS	-193	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31778533	2+3-	20	31778513	2+3-	INS	-240	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31787708	2+2-	20	31787659	2+2-	INS	-108	37	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31806228	2+2-	20	31806198	2+2-	INS	-233	26	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31821040	5+2-	20	31821082	5+2-	INS	-348	16	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	31824899	2+2-	20	31824873	2+2-	INS	-376	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31826471	3+2-	20	31826476	3+2-	INS	-109	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31829317	2+3-	20	31829333	0+2-	INS	-333	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31855811	2+2-	20	31855757	2+2-	INS	-403	32	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31858204	2+3-	20	31858155	2+3-	INS	-108	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31862115	2+2-	20	31862072	2+2-	INS	-111	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31889754	2+2-	20	31889768	2+2-	INS	-98	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31893862	2+2-	20	31893831	2+2-	INS	-103	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	31899130	3+0-	20	31899158	0+3-	INS	-244	24	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	31957888	4+3-	20	31958010	4+3-	INS	-101	22	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31976858	2+2-	20	31976844	2+2-	INS	-92	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	31978922	2+4-	20	31978949	2+4-	INS	-255	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32000202	3+2-	20	32000243	1+4-	INS	-141	30	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	32022823	2+2-	20	32022838	2+2-	INS	-96	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	32023538	2+2-	20	32023592	2+2-	INS	-97	26	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32026202	2+4-	20	32026230	2+4-	INS	-208	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32031136	2+2-	20	32031096	2+2-	INS	-101	38	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32031731	3+2-	20	32031746	3+2-	INS	-238	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32036205	3+4-	20	32036275	3+4-	INS	-217	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32041231	2+2-	20	32041234	2+2-	INS	-397	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32046321	2+2-	20	32046348	2+2-	INS	-236	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	32054810	3+2-	20	32054833	3+2-	INS	-247	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32065467	2+2-	20	32065473	2+2-	INS	-109	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32068231	2+2-	20	32068206	2+2-	INS	-375	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32081707	2+2-	20	32081756	2+2-	INS	-100	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32083329	2+3-	20	32083343	2+3-	INS	-110	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	32107377	2+2-	20	32107387	2+2-	INS	-106	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32115148	2+0-	20	32115330	0+3-	INS	-153	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32116656	2+2-	20	32116640	2+2-	INS	-125	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32119423	2+2-	20	32119388	2+2-	INS	-106	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32121053	3+3-	20	32121101	3+3-	INS	-165	27	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32133552	3+4-	20	32133620	3+4-	INS	-314	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32140508	2+3-	20	32140506	2+3-	INS	-95	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32153566	3+3-	20	32153582	3+3-	INS	-111	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32169146	2+2-	20	32169154	2+2-	INS	-229	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32172931	2+6-	20	32173047	0+2-	INS	-171	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32182099	2+2-	20	32182104	2+2-	INS	-93	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32186360	2+3-	20	32186411	2+3-	INS	-98	22	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	32202334	2+3-	20	32202397	2+3-	INS	-95	21	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	32205851	2+2-	20	32205817	2+2-	INS	-100	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32213321	4+3-	20	32213359	4+3-	INS	-108	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32218092	2+0-	20	32218218	0+2-	INS	-205	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32238561	2+4-	20	32238530	2+4-	INS	-110	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32238774	3+3-	20	32238759	3+3-	INS	-111	46	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32239081	2+0-	20	32239152	0+2-	INS	-266	28	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32244762	2+2-	20	32244754	2+2-	INS	-100	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32256387	2+3-	20	32256392	2+3-	INS	-107	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32265750	2+2-	20	32265724	2+2-	INS	-108	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32279659	48+1-	20	32282885	0+46-	DEL	3304	99	45	COLO-829BL-IL|19:COLO-829-IL|26	0.85	BreakDancerMax-0.0.1r81	|q10|o20
20	32339344	3+4-	20	32339432	0+2-	INS	-148	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32367170	2+2-	20	32367146	2+2-	INS	-374	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32369484	2+2-	20	32369480	1+3-	INS	-231	31	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	32412633	2+3-	20	32412659	2+3-	INS	-107	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32423238	2+0-	20	32423320	6+2-	INS	-230	11	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32429425	2+2-	20	32429395	2+2-	INS	-379	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32462353	2+3-	20	32462362	2+3-	INS	-110	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	32487219	3+4-	20	32487279	3+4-	INS	-242	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32493845	4+3-	20	32493925	4+3-	INS	-178	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32496842	2+2-	20	32496837	2+2-	INS	-102	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32612301	2+1-	20	32612304	1+3-	INS	-205	23	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	32639347	3+0-	20	32639429	0+3-	INS	-198	25	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32653299	3+2-	20	32653292	3+2-	INS	-118	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32653623	2+2-	20	32653616	2+2-	INS	-102	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32675472	2+3-	20	32675493	2+3-	INS	-211	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32686575	3+2-	20	32686607	3+2-	INS	-215	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	32695632	2+0-	20	32695757	0+2-	INS	-201	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32705297	5+2-	20	32707924	0+34-	DEL	2421	43	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	32705534	35+1-	20	32707924	0+32-	DEL	2433	99	29	COLO-829BL-IL|12:COLO-829-IL|17	0.74	BreakDancerMax-0.0.1r81	|q10|o20
20	32723564	2+3-	20	32723569	2+3-	INS	-94	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32734622	3+3-	20	32734646	3+3-	INS	-105	39	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32738677	3+2-	20	32738649	3+2-	INS	-117	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32746491	2+3-	20	32746496	2+3-	INS	-111	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32771518	3+4-	20	32771630	3+4-	INS	-169	23	3	COLO-829_v2_74|1:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	32780346	2+2-	20	32780310	2+2-	INS	-253	28	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32793693	2+2-	20	32793692	2+2-	INS	-228	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32804096	2+0-	20	32804272	0+2-	INS	-149	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32814258	2+2-	20	32814250	2+2-	INS	-105	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32823287	2+0-	20	32823466	0+3-	INS	-150	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32844842	2+1-	20	32844943	1+3-	INS	-188	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	32875120	2+0-	20	32875316	0+2-	INS	-137	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32907094	2+2-	20	32907105	2+2-	INS	-238	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32914603	2+2-	20	32914576	2+2-	INS	-113	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32943310	3+2-	20	32943366	3+2-	INS	-213	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	32950912	6+9-	20	32950999	6+9-	INS	-96	20	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32962103	2+2-	20	32962062	2+2-	INS	-107	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32974690	2+1-	20	32974774	3+6-	INS	-269	44	5	COLO-829_v2_74|5	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	32982717	2+2-	20	32982770	2+2-	INS	-237	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32983834	2+2-	20	32983803	2+2-	INS	-242	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	32984370	2+2-	20	32984398	2+2-	INS	-98	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	32987972	2+2-	20	32987977	2+2-	INS	-99	30	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	32997874	2+2-	20	32997898	2+2-	INS	-105	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33000448	2+3-	20	33000461	2+3-	INS	-249	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33003067	2+2-	20	33003056	2+2-	INS	-101	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33008582	3+1-	20	33008712	0+3-	INS	-163	25	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	33039368	2+2-	20	33039399	2+2-	INS	-93	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33042193	5+2-	20	33042204	1+4-	INS	-279	46	5	COLO-829_v2_74|5	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	33051304	3+1-	20	33051415	0+2-	INS	-273	27	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33062412	4+3-	20	33062449	4+3-	INS	-106	38	3	COLO-829-IL|3	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33065606	2+1-	20	33066757	0+2-	DEL	1144	39	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	33071136	3+3-	20	33071081	3+3-	INS	-309	52	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33080257	2+2-	20	33080273	2+2-	INS	-102	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33085071	5+0-	20	33085578	2+39-	DEL	323	99	5	COLO-829_v2_74|5	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	33085337	41+0-	20	33085578	2+34-	DEL	330	99	34	COLO-829BL-IL|15:COLO-829-IL|19	0.49	BreakDancerMax-0.0.1r81	|q10|o20
20	33085337	7+0-	20	33085940	0+3-	DEL	325	66	3	COLO-829_v2_74|3	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	33085337	4+0-	20	33085833	0+4-	DEL	309	93	4	COLO-829_v2_74|4	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	33095218	2+2-	20	33095203	2+2-	INS	-110	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33139830	3+3-	20	33139878	3+3-	INS	-102	36	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33145095	2+2-	20	33145044	2+2-	INS	-400	30	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33155407	3+3-	20	33155478	3+3-	INS	-161	30	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33178830	3+0-	20	33178915	0+3-	INS	-245	38	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33180931	3+4-	20	33180955	3+4-	INS	-96	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33182466	2+2-	20	33182477	2+2-	INS	-234	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33199482	2+2-	20	33199449	2+2-	INS	-383	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33208535	2+3-	20	33208561	2+3-	INS	-104	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33239014	2+1-	20	33239044	1+3-	INS	-255	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33242100	2+2-	20	33242064	2+2-	INS	-386	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33252165	3+2-	20	33252195	3+2-	INS	-369	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33275494	3+2-	20	33275540	3+2-	INS	-107	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33290867	4+3-	20	33290943	4+3-	INS	-187	26	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33317729	2+2-	20	33317695	2+2-	INS	-118	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33320885	2+0-	20	33320965	0+2-	INS	-247	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33331857	2+4-	20	33331822	2+4-	INS	-100	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33345841	2+0-	20	33346038	1+2-	INS	-131	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33353068	2+3-	20	33353053	2+3-	INS	-105	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33358106	2+0-	20	33358246	0+2-	INS	-142	17	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	33384037	3+2-	20	33384005	3+2-	INS	-106	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33392075	2+0-	20	33392092	1+3-	INS	-210	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	33398747	3+3-	20	33398832	3+3-	INS	-234	15	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33403644	2+2-	20	33403692	0+2-	INS	-272	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33414040	2+0-	20	33414076	0+2-	INS	-278	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33423724	2+2-	20	33423693	2+2-	INS	-100	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33434412	2+2-	20	33434414	2+2-	INS	-104	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33438724	2+2-	20	33438699	2+2-	INS	-108	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33442990	2+2-	20	33443009	2+2-	INS	-87	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33448042	2+2-	20	33448049	2+2-	INS	-94	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33463571	2+2-	20	33463551	2+2-	INS	-108	33	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	33464596	2+2-	20	33464559	2+2-	INS	-111	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33502630	2+0-	20	33502666	1+2-	INS	-270	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33508273	2+2-	20	33508260	2+2-	INS	-117	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33514089	2+3-	20	33514080	2+3-	INS	-120	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33530034	2+0-	20	33530129	0+2-	INS	-222	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33540935	3+2-	20	33540888	3+2-	INS	-121	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33541997	2+3-	20	33542007	2+3-	INS	-232	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33577343	2+0-	20	33577341	0+3-	INS	-239	13	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33591337	3+0-	20	33591458	3+3-	INS	-176	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33597873	2+2-	20	33597883	2+2-	INS	-103	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33598907	3+3-	20	33598893	3+3-	INS	-292	34	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	33653599	2+2-	20	33653587	2+2-	INS	-224	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33681957	2+2-	20	33681914	2+2-	INS	-112	35	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33683779	2+3-	20	33683769	2+3-	INS	-359	21	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33689344	2+0-	20	33689505	0+2-	INS	-164	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33703819	2+2-	20	33703842	2+2-	INS	-107	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33712896	2+2-	20	33712928	2+2-	INS	-90	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33716647	25+0-	20	33716930	1+28-	DEL	328	99	23	COLO-829BL-IL|12:COLO-829-IL|11	0.36	BreakDancerMax-0.0.1r81	|q10|o20
20	33716647	2+0-	20	33717249	1+3-	DEL	345	44	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	33731548	2+2-	20	33731521	2+2-	INS	-86	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33749065	2+0-	20	33749270	0+2-	INS	-117	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33752512	5+3-	20	33752592	5+3-	INS	-195	25	3	COLO-829_v2_74|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33761093	2+3-	20	33761104	2+3-	INS	-104	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33768108	2+2-	20	33768077	2+2-	INS	-123	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33778288	2+2-	20	33778297	2+2-	INS	-231	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33783983	2+2-	20	33783966	2+2-	INS	-115	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33792249	8+3-	20	33792304	8+3-	INS	-246	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33795620	2+0-	20	33795659	0+2-	INS	-266	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33825501	5+4-	20	33825624	5+4-	INS	-100	17	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33849687	2+2-	20	33849657	2+2-	INS	-105	31	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	33851575	10+2-	20	33851653	10+2-	INS	-228	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33870253	2+2-	20	33870224	2+2-	INS	-110	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33878586	3+2-	20	33878574	3+2-	INS	-116	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33880325	2+2-	20	33880446	0+2-	INS	-167	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33892591	3+0-	20	33892672	0+2-	INS	-236	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	33902651	2+2-	20	33902672	2+2-	INS	-99	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33905959	2+3-	20	33905942	2+3-	INS	-106	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33944929	2+2-	20	33944941	2+2-	INS	-245	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	33948888	3+2-	20	33948920	3+2-	INS	-241	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	33957070	2+3-	20	33957045	2+3-	INS	-391	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33982165	2+2-	20	33982132	2+2-	INS	-121	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	33985278	2+1-	20	33985348	0+2-	INS	-247	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	33989673	2+4-	20	33989727	2+4-	INS	-97	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	33995721	2+3-	20	33995722	2+3-	INS	-109	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34001696	2+2-	20	34001715	2+2-	INS	-236	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34015117	2+2-	20	34015118	2+2-	INS	-227	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34121281	5+4-	20	34121402	5+4-	INS	-173	21	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34133933	2+4-	20	34133965	2+4-	INS	-214	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34145404	2+2-	20	34145375	2+2-	INS	-241	26	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	34170471	4+2-	20	34170532	2+3-	INS	-159	33	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	34209448	2+2-	20	34209400	2+2-	INS	-109	40	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34209612	2+0-	20	34209727	0+3-	INS	-184	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34227228	2+2-	20	34227183	2+2-	INS	-106	39	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	34234286	2+2-	20	34234260	2+2-	INS	-376	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34249597	2+2-	20	34249581	2+2-	INS	-88	33	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34292494	2+2-	20	34292517	2+2-	INS	-208	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34302431	2+3-	20	34302442	2+3-	INS	-105	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34320175	2+0-	20	34320373	0+2-	INS	-120	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34336804	3+3-	20	34336801	3+3-	INS	-114	41	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34338455	2+2-	20	34338443	2+2-	INS	-249	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	34342765	2+2-	20	34342739	2+2-	INS	-96	35	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34353579	2+2-	20	34353596	2+2-	INS	-109	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34438708	2+2-	20	34438761	2+2-	INS	-333	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34458096	30+33-	20	34458348	30+33-	INS	-109	99	20	COLO-829BL-IL|7:COLO-829_v2_74|1:COLO-829-IL|12	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	34465705	2+2-	20	34465690	2+2-	INS	-114	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34475624	2+3-	20	34475643	2+3-	INS	-106	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34478356	3+0-	20	34478488	0+3-	INS	-185	33	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34522224	2+2-	20	34522182	2+2-	INS	-108	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34537564	2+2-	20	34537589	2+2-	INS	-237	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34542740	2+2-	20	34542727	2+2-	INS	-106	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34543509	3+3-	20	34543492	3+3-	INS	-95	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34569555	2+2-	20	34569555	2+2-	INS	-113	27	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34580523	3+2-	20	34580514	3+2-	INS	-119	28	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	34582233	2+2-	20	34582236	2+2-	INS	-96	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	34598374	2+2-	20	34598322	2+2-	INS	-401	31	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	34609292	3+3-	20	34609348	3+3-	INS	-186	26	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	34612980	4+3-	20	34613060	4+3-	INS	-110	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34632885	3+2-	20	34632868	3+2-	INS	-260	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	34640290	2+4-	20	34640348	2+4-	INS	-102	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34647201	2+2-	20	34647168	2+2-	INS	-117	32	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	34647726	2+1-	20	34647746	0+2-	INS	-297	19	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	34650148	2+2-	20	34650136	2+2-	INS	-234	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34658668	3+2-	20	34658689	3+2-	INS	-249	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34659207	2+3-	20	34659251	2+3-	INS	-105	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34660200	2+2-	20	34660204	2+2-	INS	-97	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34664867	2+4-	20	34664908	2+4-	INS	-107	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34665261	2+3-	20	34665227	2+3-	INS	-106	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	34665483	2+2-	20	34665448	2+2-	INS	-109	32	2	COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	34671502	2+0-	20	34671666	1+2-	INS	-169	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34678023	5+4-	20	34678128	5+4-	INS	-199	22	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34682783	2+2-	20	34682814	2+2-	INS	-248	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34685830	3+0-	20	34685985	1+4-	INS	-154	47	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34693289	2+2-	20	34693272	2+2-	INS	-107	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	34698844	5+3-	20	34698872	5+3-	INS	-368	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34734242	3+1-	20	34734306	0+2-	INS	-268	25	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	34759520	2+1-	20	34759625	2+6-	INS	-121	13	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34769159	2+3-	20	34769188	2+3-	INS	-230	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34775209	4+4-	20	34775257	4+4-	INS	-243	36	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34775833	2+2-	20	34775843	2+2-	INS	-103	26	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	34785116	3+3-	20	34785155	3+3-	INS	-111	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	34794315	2+2-	20	34794306	2+2-	INS	-108	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34802172	3+2-	20	34802155	3+2-	INS	-111	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34830213	2+2-	20	34830254	2+2-	INS	-198	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34863165	2+2-	20	34863161	2+2-	INS	-115	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34893959	2+1-	20	34893989	0+2-	INS	-256	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34909149	2+2-	20	34909154	2+2-	INS	-86	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34913381	2+2-	20	34913344	2+2-	INS	-387	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34917802	2+3-	20	34917844	2+3-	INS	-100	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34920141	4+1-	20	34920291	0+4-	DEL	105	69	3	COLO-829BL-IL|2:COLO-829-IL|1	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	34935671	2+2-	20	34935627	2+2-	INS	-112	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	34939027	2+0-	20	34939085	1+2-	INS	-280	29	2	COLO-829_v2_74|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	34943793	2+2-	20	34943757	2+2-	INS	-386	25	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	34952114	18+2-	20	34952173	18+2-	INS	-216	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34954175	2+3-	20	34954133	2+3-	INS	-111	34	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	34979078	2+2-	20	34979090	2+2-	INS	-110	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	34982158	1+3-	20	34982496	1+3-	INV	241	53	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35009088	4+0-	20	35009092	10+13-	INS	-95	53	6	COLO-829BL-IL|2:COLO-829-IL|4	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	35027421	2+12-	20	35042567	0+11-	INV	15096	99	11	COLO-829BL-IL|3:COLO-829-IL|8	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	35028016	4+0-	20	35041288	5+1-	INV	13247	99	4	COLO-829BL-IL|1:COLO-829-IL|3	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	35028877	1+3-	20	35034557	1+3-	INV	5607	50	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	35039547	4+7-	20	35039602	4+7-	INS	-94	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35045701	2+4-	20	35045757	2+4-	INS	-111	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35062902	2+1-	20	35063000	0+4-	DEL	92	46	2	COLO-829BL-IL|2	0.40	BreakDancerMax-0.0.1r81	|q10|o20
20	35083595	4+5-	20	35083636	4+5-	INS	-367	39	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35098016	2+1-	20	35098429	3+3-	DEL	77	49	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	35101978	3+0-	20	35101968	1+3-	INS	-234	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	35105989	2+2-	20	35105949	2+2-	INS	-106	34	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35111196	2+0-	20	35111313	0+2-	INS	-194	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35115275	2+2-	20	35115255	2+2-	INS	-370	22	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	35148635	2+2-	20	35148679	2+2-	INS	-94	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35157177	2+0-	20	35157199	0+2-	INS	-296	20	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	35158776	2+0-	20	35158786	0+2-	INS	-292	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35175122	4+1-	20	35175166	1+4-	INS	-237	37	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	35177652	2+2-	20	35177674	2+2-	INS	-97	24	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35192543	2+3-	20	35192527	2+3-	INS	-101	33	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35216740	2+2-	20	35216777	2+2-	INS	-233	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35226901	2+2-	20	35226887	2+2-	INS	-111	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35235231	2+2-	20	35235253	2+2-	INS	-94	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35239470	4+3-	20	35239504	4+3-	INS	-100	38	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35245496	2+2-	20	35245493	2+2-	INS	-96	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35249072	50+0-	20	35249518	0+3-	DEL	310	42	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	35249072	48+0-	20	35249332	0+47-	DEL	319	99	47	COLO-829BL-IL|14:COLO-829-IL|33	0.48	BreakDancerMax-0.0.1r81	|q10|o20
20	35253948	2+0-	20	35253989	0+2-	INS	-295	27	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35258671	2+3-	20	35258711	2+3-	INS	-213	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35264676	2+2-	20	35264620	2+2-	INS	-117	40	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35279163	2+3-	20	35279166	2+3-	INS	-95	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35280965	2+3-	20	35280980	2+3-	INS	-225	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35288780	2+2-	20	35288803	2+2-	INS	-361	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35298849	2+3-	20	35298890	2+3-	INS	-89	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	35301170	2+2-	20	35301184	2+2-	INS	-102	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35303834	2+2-	20	35303855	0+2-	INS	-292	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35313291	2+2-	20	35313253	2+2-	INS	-98	37	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35316884	3+2-	20	35316930	3+2-	INS	-100	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35345026	2+3-	20	35345069	2+3-	INS	-198	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35345501	2+2-	20	35345487	2+2-	INS	-107	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35354904	2+2-	20	35354879	2+2-	INS	-108	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35356353	3+1-	20	35356474	0+2-	INS	-187	42	3	COLO-829_v2_74|2:COLO-829-IL|1	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	35357678	4+3-	20	35357759	4+3-	INS	-204	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35385198	2+2-	20	35385163	2+2-	INS	-113	32	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	35401961	2+2-	20	35401954	2+2-	INS	-100	32	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35405368	2+3-	20	35405374	2+3-	INS	-112	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	35406012	2+2-	20	35405961	2+2-	INS	-255	32	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	35407176	2+0-	20	35407316	0+2-	INS	-184	22	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	35423663	11+1-	20	35423670	0+10-	DEL	100	99	10	COLO-829BL-IL|5:COLO-829-IL|5	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	35437381	3+3-	20	35437470	3+3-	INS	-111	18	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35461056	3+3-	20	35461093	3+3-	INS	-216	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35462025	2+2-	20	35462024	2+2-	INS	-231	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35523395	2+3-	20	35523420	2+3-	INS	-107	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35542975	3+0-	20	35543035	0+3-	INS	-235	30	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	35550555	4+3-	20	35550627	0+2-	INS	-136	22	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35555458	2+2-	20	35555519	1+3-	INS	-175	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35555769	2+0-	20	35555863	0+2-	INS	-223	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35559814	3+3-	20	35559823	3+3-	INS	-93	39	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35563625	3+1-	20	35563688	0+3-	INS	-256	34	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35565682	4+1-	20	35565668	0+4-	INS	-257	35	4	COLO-829_v2_74|3:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	35572871	3+1-	20	35573037	1+2-	INS	-127	27	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35576298	2+2-	20	35576288	2+2-	INS	-242	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35641281	3+2-	20	35641339	3+2-	INS	-97	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35647481	2+2-	20	35647481	2+2-	INS	-250	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35654292	3+1-	20	35654304	0+3-	INS	-297	29	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35655078	2+0-	20	35655099	2+4-	INS	-262	20	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35663447	2+2-	20	35663416	2+2-	INS	-102	32	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	35672819	5+7-	20	35672907	5+7-	ITX	-129	34	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35674826	3+2-	20	35674821	3+2-	INS	-92	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35683848	2+1-	20	35683865	1+3-	INS	-256	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35697170	3+3-	20	35697199	3+3-	INS	-262	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35697485	2+2-	20	35697443	2+2-	INS	-392	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35720406	3+4-	20	35720445	3+4-	INS	-280	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	35721380	2+4-	20	35721422	2+4-	INS	-100	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35744012	3+3-	20	35744022	3+3-	INS	-285	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	35747094	2+2-	20	35747106	2+2-	INS	-213	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35747244	3+2-	20	35747261	3+2-	INS	-110	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	35786887	2+2-	20	35786843	2+2-	INS	-113	35	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	35795428	4+2-	20	35795396	4+2-	INS	-250	27	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35799372	2+2-	20	35799351	2+2-	INS	-371	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35834934	2+2-	20	35834974	2+2-	INS	-87	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	35869264	2+2-	20	35869263	2+2-	INS	-97	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35885582	2+2-	20	35885546	2+2-	INS	-239	28	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	35924432	3+1-	20	35924448	0+2-	INS	-240	33	3	COLO-829_v2_74|2:COLO-829-IL|1	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	35936593	2+0-	20	35936637	0+2-	INS	-273	20	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	35950143	2+2-	20	35950093	2+2-	INS	-118	37	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	35955536	13+5-	20	35955638	13+5-	INS	-101	18	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35976217	3+0-	20	35976295	0+3-	INS	-230	30	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35987029	3+1-	20	35987211	0+2-	INS	-125	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	35996733	2+2-	20	35996731	2+2-	INS	-248	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36001279	2+2-	20	36001254	2+2-	INS	-89	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36005271	2+3-	20	36005304	2+3-	INS	-99	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36020702	2+2-	20	36020668	2+2-	INS	-100	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36021470	2+2-	20	36021460	2+2-	INS	-90	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36023088	3+0-	20	36023164	0+4-	INS	-246	31	3	COLO-829_v2_74|3	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	36052271	2+2-	20	36052256	2+2-	INS	-384	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36057106	2+1-	20	36057236	0+2-	INS	-198	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36074176	2+2-	20	36074176	2+2-	INS	-91	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36080005	2+2-	20	36079979	2+2-	INS	-101	35	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36086652	2+3-	20	36086691	2+3-	INS	-113	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36093281	2+3-	20	36093317	2+3-	INS	-373	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36099842	2+4-	20	36099849	2+4-	INS	-100	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36124342	4+3-	20	36124376	4+3-	INS	-191	28	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36132077	2+3-	20	36132124	2+3-	INS	-102	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36159467	2+3-	20	36159438	2+3-	INS	-378	24	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36189633	2+2-	20	36189619	2+2-	INS	-108	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36202040	2+0-	20	36202140	0+2-	INS	-232	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36208415	2+2-	20	36208385	2+2-	INS	-105	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36217240	2+2-	20	36217238	2+2-	INS	-237	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36234158	2+2-	20	36234097	2+2-	INS	-411	36	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36242768	2+2-	20	36242777	2+2-	INS	-112	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36246087	3+2-	20	36246176	1+2-	INS	-224	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36256189	34+41-	20	36256595	34+41-	INS	-99	55	7	COLO-829BL-IL|3:COLO-829-IL|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36258673	3+2-	20	36258731	3+2-	INS	-347	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36282919	2+1-	20	36282904	1+2-	INS	-346	19	2	COLO-829_v2_74|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	36309547	2+2-	20	36309495	2+2-	INS	-401	31	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36336719	3+1-	20	36336931	0+2-	INS	-105	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36338844	2+2-	20	36338879	2+2-	INS	-94	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36349788	2+2-	20	36349764	2+2-	INS	-93	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36365339	2+2-	20	36365314	2+2-	INS	-113	34	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36370533	2+2-	20	36370588	2+2-	INS	-103	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36375973	8+1-	20	36376046	14+21-	ITX	-144	99	10	COLO-829BL-IL|5:COLO-829-IL|5	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	36376676	3+1-	20	36376755	0+2-	INS	-315	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36386110	3+1-	20	36386196	1+3-	INS	-178	48	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36400996	2+2-	20	36400964	2+2-	INS	-243	27	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36404533	2+3-	20	36404477	2+3-	INS	-120	38	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36411182	2+0-	20	36411226	0+2-	INS	-278	21	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36425073	2+2-	20	36425022	2+2-	INS	-110	36	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36431574	3+0-	20	36431671	0+3-	INS	-191	22	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36449449	3+2-	20	36449505	3+2-	INS	-88	26	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36452540	3+3-	20	36452598	3+3-	INS	-239	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36462554	2+3-	20	36462533	2+3-	INS	-103	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36475586	2+2-	20	36475528	2+2-	INS	-115	45	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36510412	2+2-	20	36510359	2+2-	INS	-403	31	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36519527	2+2-	20	36519549	2+2-	INS	-106	24	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36520588	3+4-	20	36520628	3+4-	INS	-204	28	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36525684	2+0-	20	36525914	0+2-	DEL	187	45	2	COLO-829BL-IL|1:COLO-829-IL|1	0.22	BreakDancerMax-0.0.1r81	|q10|o20
20	36537525	3+3-	20	36537565	3+3-	INS	-224	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36541965	2+4-	20	36541945	2+4-	INS	-85	33	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36548494	2+2-	20	36548447	2+2-	INS	-105	40	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36553956	2+2-	20	36553955	2+2-	INS	-89	31	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36560274	2+5-	20	36560270	2+5-	INS	-93	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36581695	2+2-	20	36581687	2+2-	INS	-93	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36584192	2+3-	20	36584204	2+3-	INS	-222	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36622486	2+2-	20	36622497	2+2-	INS	-231	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36642515	2+2-	20	36642499	2+2-	INS	-410	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36648880	2+0-	20	36648875	0+2-	INS	-308	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36670750	2+3-	20	36670729	2+3-	INS	-248	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36682011	2+3-	20	36681999	2+3-	INS	-103	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36685977	3+4-	20	36686014	3+4-	INS	-275	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36688385	2+3-	20	36688395	2+3-	INS	-233	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36689415	18+20-	20	36689682	18+20-	DEL	91	99	15	COLO-829BL-IL|5:COLO-829-IL|10	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36693452	3+2-	20	36693454	3+2-	INS	-99	26	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36714268	2+0-	20	36714291	0+2-	INS	-291	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36715412	59+48-	20	36715414	0+2-	INS	-220	99	36	COLO-829BL-IL|2:COLO-829_v2_74|27:COLO-829-IL|7	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	36715656	3+5-	20	36715721	3+5-	INS	-204	25	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36722423	3+1-	20	36722514	0+2-	INS	-175	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36733237	4+2-	20	36733243	1+3-	INS	-211	43	5	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	36777752	2+3-	20	36777744	2+3-	INS	-250	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36813150	2+2-	20	36813270	1+2-	INS	-150	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36831523	2+3-	20	36831520	2+3-	INS	-251	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36831861	3+1-	20	36831910	1+3-	INS	-186	40	4	COLO-829_v2_74|2:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36849005	2+3-	20	36849029	2+3-	INS	-112	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36860356	2+2-	20	36860331	2+2-	INS	-100	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36877046	3+3-	20	36877185	1+3-	INS	-181	18	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36912029	2+2-	20	36911997	2+2-	INS	-235	27	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36915447	3+0-	20	36915468	0+3-	INS	-300	34	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36939943	2+3-	20	36940007	2+3-	INS	-202	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36942676	3+2-	20	36942725	3+2-	INS	-243	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36944113	3+3-	20	36944112	3+3-	INS	-200	35	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36948817	2+2-	20	36948841	2+2-	INS	-243	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	36950537	2+0-	20	36950671	1+3-	INS	-141	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36954580	2+2-	20	36954566	2+2-	INS	-108	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	36957866	4+4-	20	36957924	4+4-	INS	-98	35	3	COLO-829BL-IL|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	36965579	6+6-	20	36965605	6+6-	INS	-95	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36971981	2+2-	20	36971964	2+2-	INS	-367	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	36986624	2+0-	20	36986698	2+3-	INS	-200	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	37002483	2+0-	20	37002698	0+2-	INS	-119	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37022920	2+2-	20	37022917	2+2-	INS	-231	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37032026	4+3-	20	37032148	4+3-	INS	-331	12	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37054591	3+0-	20	37054605	0+3-	INS	-294	31	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37064887	2+2-	20	37064861	2+2-	INS	-104	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37072688	2+0-	20	37072716	2+4-	INS	-229	32	4	COLO-829_v2_74|3:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	37095478	2+2-	20	37095469	2+2-	INS	-108	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37137266	3+2-	20	37137233	3+2-	INS	-107	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37143268	2+0-	20	37143299	0+2-	INS	-269	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37153839	2+2-	20	37153827	2+2-	INS	-100	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37155700	3+1-	20	37155708	1+2-	INS	-241	14	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37190514	3+2-	20	37190540	0+2-	INS	-234	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37191024	2+0-	20	37191197	0+2-	INS	-150	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37193240	2+2-	20	37193219	2+2-	INS	-371	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37202462	3+3-	20	37202512	3+3-	INS	-285	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37214540	3+1-	20	37214543	0+2-	INS	-246	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37227259	2+2-	20	37227268	2+2-	INS	-92	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37240382	2+0-	20	37240399	1+2-	INS	-254	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37249037	2+3-	20	37249039	2+3-	INS	-100	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37260544	2+2-	20	37260515	2+2-	INS	-103	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37284767	3+0-	20	37284791	0+3-	INS	-295	35	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37301182	2+2-	20	37301213	2+2-	INS	-243	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37309898	2+2-	20	37309906	2+2-	INS	-373	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37315194	3+2-	20	37315161	3+2-	INS	-243	25	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37327772	3+0-	20	37327926	0+3-	INS	-168	37	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37329225	2+2-	20	37329239	2+2-	INS	-92	29	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37339552	2+0-	20	37339682	1+3-	INS	-125	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37356871	2+2-	20	37356874	2+2-	INS	-99	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37360434	3+5-	20	37360542	3+5-	INS	-92	32	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37388162	4+4-	20	37388174	4+4-	INS	-88	55	4	COLO-829BL-IL|2:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37400588	9+1-	20	37400865	1+30-	DEL	85	99	9	COLO-829_v2_74|9	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	37400850	21+0-	20	37400865	0+20-	DEL	93	99	20	COLO-829BL-IL|9:COLO-829-IL|11	0.19	BreakDancerMax-0.0.1r81	|q10|o20
20	37419844	4+3-	20	37419876	4+3-	INS	-287	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37435830	2+3-	20	37435798	2+3-	INS	-106	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37458464	2+2-	20	37458448	2+2-	INS	-229	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37511887	2+2-	20	37511882	2+2-	INS	-242	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37512572	4+3-	20	37512592	4+3-	INS	-111	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37515613	2+0-	20	37515763	1+3-	INS	-113	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37528999	2+2-	20	37529040	2+2-	INS	-350	16	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37549821	3+3-	20	37549863	3+3-	INS	-110	37	3	COLO-829-IL|3	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37550714	2+3-	20	37550747	2+3-	INS	-101	23	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37578072	2+2-	20	37578041	2+2-	INS	-381	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37616764	2+2-	20	37616807	2+2-	INS	-223	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37630413	2+2-	20	37630443	2+2-	INS	-85	28	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37651559	2+2-	20	37651546	2+2-	INS	-377	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37663614	2+3-	20	37663618	2+3-	INS	-105	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37678004	2+2-	20	37677961	2+2-	INS	-109	39	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37680702	3+3-	20	37680700	3+3-	INS	-98	41	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37700946	2+0-	20	37701020	0+2-	INS	-254	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37705264	2+3-	20	37705300	2+3-	INS	-99	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37720567	3+3-	20	37720623	3+3-	INS	-107	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37727637	2+2-	20	37727612	2+2-	INS	-115	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37753295	2+3-	20	37753328	2+3-	INS	-245	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37758209	2+0-	20	37758343	0+2-	INS	-170	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37770809	2+0-	20	37771178	1+39-	DEL	133	46	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37771098	39+0-	20	37771178	1+37-	DEL	135	99	35	COLO-829BL-IL|11:COLO-829-IL|24	0.28	BreakDancerMax-0.0.1r81	|q10|o20
20	37771098	4+0-	20	37771465	0+4-	DEL	147	65	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	37776111	3+3-	20	37776100	3+3-	INS	-96	44	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37811177	3+1-	20	37811276	0+2-	INS	-164	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37817474	3+2-	20	37817499	1+3-	INS	-241	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	37824281	2+2-	20	37824260	2+2-	INS	-102	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37825728	2+0-	20	37825843	0+3-	INS	-201	21	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	37834071	2+2-	20	37834019	2+2-	INS	-114	38	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37850526	2+3-	20	37850540	2+3-	INS	-99	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37851225	2+2-	20	37851190	2+2-	INS	-108	36	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37886730	3+1-	20	37886827	1+4-	INS	-214	29	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37887638	2+2-	20	37887652	2+2-	INS	-219	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	37888029	2+0-	20	37888115	0+2-	INS	-229	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37897794	2+2-	20	37897782	2+2-	INS	-101	32	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37901340	2+0-	20	37901492	0+2-	INS	-171	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37919750	2+3-	20	37919778	2+3-	INS	-99	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37928676	2+2-	20	37928622	2+2-	INS	-110	37	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37933271	2+2-	20	37933285	2+2-	INS	-103	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37937695	2+2-	20	37937668	2+2-	INS	-259	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37939311	3+2-	20	37939319	3+2-	INS	-111	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37946540	23+12-	20	37946632	1+12-	INS	-105	99	12	COLO-829BL-IL|4:COLO-829-IL|8	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	37953614	2+2-	20	37953607	2+2-	INS	-234	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	37964877	3+2-	20	37964921	3+2-	INS	-92	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	37985208	3+2-	20	37985269	3+2-	INS	-107	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38014928	3+2-	20	38014905	3+2-	INS	-243	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38015074	2+3-	20	38015083	2+3-	INS	-241	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38026427	2+1-	20	38026465	1+2-	INS	-299	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38034897	2+2-	20	38034873	2+2-	INS	-115	30	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	38049182	2+2-	20	38049207	2+2-	INS	-255	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38059995	2+2-	20	38060029	2+2-	INS	-92	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38085746	3+3-	20	38085727	1+4-	INS	-285	28	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38106247	4+4-	20	38106268	4+4-	INS	-259	42	4	COLO-829_v2_74|2:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38117995	3+2-	20	38118217	1+3-	INS	-116	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	38120106	2+2-	20	38120060	2+2-	INS	-104	40	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	38127826	2+0-	20	38127903	0+2-	INS	-264	31	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38161675	3+2-	20	38161672	3+2-	INS	-107	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38171316	2+2-	20	38171337	2+2-	INS	-92	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38178245	2+2-	20	38178223	2+2-	INS	-97	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	38178809	3+2-	20	38178788	3+2-	INS	-89	34	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38180883	2+0-	20	38180908	1+3-	INS	-207	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38181962	2+2-	20	38181997	2+2-	INS	-93	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38192835	2+2-	20	38192815	2+2-	INS	-369	22	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	38195151	3+1-	20	38195149	1+3-	INS	-207	35	4	COLO-829_v2_74|2:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	38202878	3+2-	20	38202929	1+3-	INS	-177	45	4	COLO-829_v2_74|2:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	38220175	2+2-	20	38220129	2+2-	INS	-396	28	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	38224230	3+0-	20	38224386	1+3-	INS	-150	33	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	38231744	3+3-	20	38231781	3+3-	INS	-188	28	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38238471	4+3-	20	38238495	4+3-	INS	-190	35	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38249830	2+1-	20	38249932	0+3-	INS	-220	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38262681	3+3-	20	38262745	3+3-	INS	-104	35	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38266072	3+2-	20	38266073	3+2-	INS	-109	31	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38284163	2+0-	20	38284145	0+2-	INS	-234	30	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38286163	2+0-	20	38286240	0+2-	INS	-226	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38297343	2+2-	20	38297312	2+2-	INS	-112	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38157219	4+0-	20	38332965	0+6-	DEL	175726	70	4	COLO-829BL-IL|2:COLO-829-IL|2	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	38330657	3+3-	20	38330710	3+3-	INS	-92	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38340921	3+1-	20	38341074	0+3-	INS	-163	29	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38363789	2+2-	20	38363771	2+2-	INS	-100	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38365912	2+2-	20	38365889	2+2-	INS	-372	23	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	38368386	2+0-	20	38368389	0+2-	INS	-320	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38372072	2+2-	20	38372106	2+2-	INS	-99	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38385443	3+3-	20	38385487	3+3-	INS	-111	37	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38396658	2+3-	20	38396646	2+3-	INS	-98	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38401345	2+2-	20	38401324	2+2-	INS	-110	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38418725	2+2-	20	38418702	2+2-	INS	-372	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38419605	4+1-	20	38419650	0+2-	INS	-213	27	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38425655	2+3-	20	38425721	2+3-	INS	-230	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	38437390	3+3-	20	38437363	3+3-	INS	-93	46	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38460304	2+2-	20	38460276	2+2-	INS	-378	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38461120	2+1-	20	38461166	0+2-	INS	-267	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38465438	2+3-	20	38465450	2+3-	INS	-113	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38473531	3+1-	20	38473616	0+2-	INS	-168	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38484586	3+4-	20	38484684	3+4-	INS	-223	15	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	38493870	2+2-	20	38493845	2+2-	INS	-94	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38509122	2+2-	20	38509081	2+2-	INS	-110	34	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	38513764	2+2-	20	38513734	2+2-	INS	-105	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38518414	2+2-	20	38518378	2+2-	INS	-93	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38521990	2+0-	20	38522073	12+7-	INS	-194	13	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	38536290	2+2-	20	38536321	2+2-	INS	-90	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38569241	3+0-	20	38569224	0+4-	INS	-295	26	3	COLO-829_v2_74|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	38574146	3+3-	20	38574209	3+3-	INS	-104	35	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38575542	3+2-	20	38575546	3+2-	INS	-125	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38577637	2+2-	20	38577616	2+2-	INS	-250	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38594448	3+3-	20	38594453	3+3-	INS	-265	32	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38599559	3+0-	20	38599656	0+3-	INS	-186	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38600614	3+3-	20	38600670	0+2-	INS	-218	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38605948	3+3-	20	38606021	0+2-	INS	-160	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38639611	2+0-	20	38639659	0+2-	INS	-259	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38651563	3+0-	20	38651554	1+4-	INS	-239	38	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	38658008	3+4-	20	38658002	3+4-	INS	-196	36	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38660464	4+2-	20	38660460	4+2-	INS	-108	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38665969	2+2-	20	38665942	2+2-	INS	-377	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38668229	3+2-	20	38668221	1+2-	INS	-300	22	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38690095	3+2-	20	38690058	3+2-	INS	-392	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38696698	4+1-	20	38696783	1+3-	INS	-242	35	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38705881	2+2-	20	38705847	2+2-	INS	-118	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	38727870	2+1-	20	38727863	1+3-	INS	-249	35	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	38744803	2+2-	20	38744781	2+2-	INS	-234	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38748220	2+0-	20	38748368	0+2-	INS	-179	23	2	COLO-829_v2_74|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	38763733	3+0-	20	38763755	0+3-	INS	-305	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38771028	2+2-	20	38770988	2+2-	INS	-390	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38771578	5+3-	20	38771604	5+3-	INS	-279	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38781649	2+3-	20	38781688	2+3-	INS	-245	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38788042	3+2-	20	38788057	0+2-	INS	-184	23	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38790637	3+3-	20	38790694	3+3-	INS	-106	35	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38815985	2+2-	20	38815956	2+2-	INS	-99	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38828344	2+0-	20	38828401	1+3-	INS	-175	30	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38835944	2+2-	20	38835949	2+2-	INS	-229	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38837877	2+3-	20	38837870	2+3-	INS	-239	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38843077	2+2-	20	38843069	2+2-	INS	-89	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	38893262	3+3-	20	38893348	3+3-	INS	-273	21	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38910077	2+0-	20	38910170	1+2-	INS	-209	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38910420	2+3-	20	38910405	2+3-	INS	-107	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	38913428	3+2-	20	38913447	3+2-	INS	-376	18	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	38915789	2+2-	20	38915765	2+2-	INS	-113	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38927987	2+2-	20	38927958	2+2-	INS	-106	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38931248	2+0-	20	38931303	0+2-	INS	-267	21	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	38964616	2+0-	20	38964820	0+2-	INS	-125	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38984335	4+0-	20	38984351	0+2-	INS	-247	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	38994943	2+2-	20	38994892	2+2-	INS	-257	30	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39005046	3+0-	20	39005147	1+5-	INS	-187	36	4	COLO-829_v2_74|3:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	39007352	2+2-	20	39007385	2+2-	INS	-206	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39007565	2+2-	20	39007648	2+2-	INS	-98	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39011112	3+2-	20	39011104	0+2-	INS	-206	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39015851	3+1-	20	39015909	0+2-	INS	-153	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39025691	2+0-	20	39025914	0+2-	INS	-116	29	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39030021	2+2-	20	39030042	2+2-	INS	-107	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39041715	2+2-	20	39041683	2+2-	INS	-120	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39045006	2+2-	20	39044996	2+2-	INS	-116	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39052866	2+0-	20	39052917	0+2-	INS	-270	21	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	39061314	2+2-	20	39061338	2+2-	INS	-101	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39084794	4+3-	20	39084850	4+3-	INS	-95	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39085337	4+2-	20	39085348	4+2-	INS	-222	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39092280	2+2-	20	39092248	2+2-	INS	-99	36	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39102035	3+4-	20	39102128	3+4-	INS	-157	24	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39112641	6+5-	20	39112759	0+3-	INS	-226	25	4	COLO-829_v2_74|3:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39116573	3+2-	20	39116578	3+2-	INS	-101	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39143508	2+2-	20	39143523	2+2-	INS	-241	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39150805	2+2-	20	39150769	2+2-	INS	-386	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39163455	2+2-	20	39163462	2+2-	INS	-251	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39172627	2+3-	20	39172632	2+3-	INS	-228	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39195778	2+2-	20	39195785	2+2-	INS	-104	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39207890	3+2-	20	39207938	2+3-	INS	-145	24	3	COLO-829_v2_74|1:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	39220237	3+3-	20	39220268	3+3-	INS	-356	28	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39221194	2+0-	20	39221260	1+3-	INS	-189	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	39229381	2+2-	20	39229474	1+3-	INS	-254	25	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39255029	2+2-	20	39255006	2+2-	INS	-108	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39257772	3+3-	20	39257787	3+3-	INS	-110	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39262830	2+2-	20	39262796	2+2-	INS	-97	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39263770	2+0-	20	39263956	2+3-	INS	-116	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39275809	2+2-	20	39275799	2+2-	INS	-105	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39280754	8+2-	20	39280907	8+2-	INS	-95	17	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39284974	3+2-	20	39284967	3+2-	INS	-113	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39287037	3+3-	20	39287122	3+3-	INS	-89	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39289842	2+2-	20	39289828	2+2-	INS	-104	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	39303110	2+1-	20	39303156	0+2-	INS	-262	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39304864	2+3-	20	39304840	2+3-	INS	-238	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39306535	2+0-	20	39306626	2+5-	INS	-156	24	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	39306643	3+1-	20	39306626	1+2-	INS	-323	22	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	39318672	2+0-	20	39318815	1+2-	INS	-150	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39319169	2+3-	20	39319207	2+3-	INS	-242	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39320743	2+1-	20	39320756	1+3-	INS	-190	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	39329422	3+0-	20	39329467	1+4-	INS	-222	43	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	39340646	3+3-	20	39340685	3+3-	INS	-232	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39349672	2+0-	20	39349847	0+2-	INS	-143	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39364463	2+2-	20	39364468	2+2-	INS	-248	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39373969	2+0-	20	39374006	0+3-	INS	-269	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39391085	3+2-	20	39391063	3+2-	INS	-254	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39398688	2+5-	20	39398757	2+5-	INS	-100	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39414684	2+2-	20	39414670	2+2-	INS	-102	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39427634	2+2-	20	39427614	2+2-	INS	-370	22	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39434339	2+3-	20	39434323	2+3-	INS	-92	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39441298	2+4-	20	39441293	2+4-	INS	-109	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39456076	2+0-	20	39456194	0+2-	INS	-186	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39474245	3+2-	20	39474251	3+2-	INS	-220	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39477935	2+2-	20	39477895	2+2-	INS	-113	34	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39490664	2+3-	20	39490677	2+3-	INS	-113	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39491653	2+2-	20	39491620	2+2-	INS	-110	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39498927	3+1-	20	39498994	0+3-	INS	-227	29	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39504727	2+1-	20	39504825	0+2-	INS	-212	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39507200	4+3-	20	39507305	4+3-	INS	-192	14	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39517530	2+3-	20	39517542	2+3-	INS	-104	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39518163	2+2-	20	39518116	2+2-	INS	-122	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39520791	2+2-	20	39520763	2+2-	INS	-93	35	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	39524241	2+1-	20	39524369	0+2-	INS	-181	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39561015	2+0-	20	39561109	0+2-	INS	-239	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39576368	2+0-	20	39576390	0+2-	INS	-288	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39577371	2+0-	20	39577362	0+2-	INS	-207	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39584479	2+3-	20	39584522	2+3-	INS	-212	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39588238	2+1-	20	39588415	0+2-	INS	-151	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39609099	2+2-	20	39609118	2+2-	INS	-91	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39617248	3+1-	20	39617334	0+3-	DEL	94	35	2	COLO-829-IL|2	0.33	BreakDancerMax-0.0.1r81	|q10|o20
20	39657140	2+2-	20	39657138	2+2-	INS	-99	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39658362	2+2-	20	39658318	2+2-	INS	-260	28	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39671608	4+0-	20	39671663	1+2-	INS	-259	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39671608	2+0-	20	39671738	3+3-	INS	-217	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39678402	2+2-	20	39678361	2+2-	INS	-105	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39693080	2+3-	20	39693172	2+3-	INS	-173	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39694615	13+20-	20	39694590	13+20-	INS	-96	99	6	COLO-829BL-IL|1:COLO-829-IL|5	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	39712536	2+1-	20	39712641	0+2-	INS	-185	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39724676	2+1-	20	39724783	0+2-	INS	-221	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39756676	5+0-	20	39756680	22+25-	INS	-124	99	25	COLO-829BL-IL|8:COLO-829_v2_74|6:COLO-829-IL|11	0.19	BreakDancerMax-0.0.1r81	|q10|o20
20	39761712	2+2-	20	39761724	2+2-	INS	-95	29	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39765424	4+3-	20	39765416	4+3-	INS	-96	44	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39766218	2+2-	20	39766219	2+2-	INS	-97	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39770787	2+2-	20	39770798	2+2-	INS	-101	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39775098	2+3-	20	39775147	2+3-	INS	-241	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39778366	2+3-	20	39778346	2+3-	INS	-106	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39780334	3+1-	20	39780387	1+2-	INS	-143	20	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39797489	2+0-	20	39797578	0+2-	INS	-223	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39822555	2+0-	20	39822607	0+3-	INS	-249	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39830893	3+3-	20	39830945	3+3-	INS	-96	42	3	COLO-829BL-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39832956	2+2-	20	39832977	2+2-	INS	-93	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39864475	5+3-	20	39864516	5+3-	INS	-103	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39895333	2+2-	20	39895297	2+2-	INS	-248	26	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	39905800	3+2-	20	39905852	3+2-	INS	-234	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39944589	3+3-	20	39944560	3+3-	INS	-113	47	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39945690	2+0-	20	39945734	0+2-	INS	-268	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39955398	2+0-	20	39955567	0+2-	INS	-133	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39964137	2+2-	20	39964142	2+2-	INS	-110	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	39978945	2+0-	20	39978936	1+4-	INS	-222	21	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	39984717	2+2-	20	39984696	2+2-	INS	-244	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	39990289	2+2-	20	39990273	2+2-	INS	-87	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40014951	2+2-	20	40014941	2+2-	INS	-93	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40039085	2+2-	20	40039052	2+2-	INS	-107	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40059774	2+2-	20	40059763	2+2-	INS	-245	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40077380	2+3-	20	40077399	2+3-	INS	-364	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40099114	2+1-	20	40099164	1+3-	INS	-227	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40107505	2+2-	20	40107555	2+2-	INS	-239	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40108998	3+0-	20	40109129	0+3-	INS	-188	33	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40118837	2+0-	20	40118881	0+3-	INS	-286	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40119860	3+2-	20	40119991	3+2-	INS	-216	11	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40161013	2+0-	20	40161067	1+2-	INS	-248	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40167074	2+3-	20	40167098	2+3-	INS	-235	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40169920	3+2-	20	40169992	3+2-	INS	-226	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40179047	2+0-	20	40179054	0+2-	INS	-325	25	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	40182620	2+2-	20	40182591	2+2-	INS	-114	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40183814	3+2-	20	40183855	3+2-	INS	-97	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40187367	2+1-	20	40187417	2+3-	INS	-176	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40187837	2+5-	20	40187955	2+5-	INS	-94	22	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40188609	2+2-	20	40188609	2+2-	INS	-93	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40202745	2+1-	20	40202841	0+2-	INS	-236	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40217209	2+0-	20	40217318	0+2-	INS	-215	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40223332	2+0-	20	40223398	2+3-	INS	-265	27	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	40224617	2+3-	20	40224667	2+3-	INS	-110	22	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40232326	2+3-	20	40232313	2+3-	INS	-363	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40241370	2+2-	20	40241386	2+2-	INS	-103	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40247775	2+2-	20	40247764	2+2-	INS	-113	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40250377	2+2-	20	40250412	2+2-	INS	-97	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40253311	2+0-	20	40253377	0+3-	INS	-215	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40254602	2+2-	20	40254635	2+2-	INS	-207	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40265729	2+2-	20	40265739	2+2-	INS	-360	18	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40277731	2+3-	20	40277797	2+3-	INS	-91	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40292621	2+2-	20	40292570	2+2-	INS	-400	30	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40292822	2+0-	20	40292880	0+2-	INS	-258	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40299772	2+3-	20	40299737	2+3-	INS	-98	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40302377	2+1-	20	40302453	0+4-	INS	-254	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40305310	3+4-	20	40305336	3+4-	INS	-261	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40305981	2+2-	20	40305983	2+2-	INS	-99	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40315892	2+2-	20	40315891	2+2-	INS	-98	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40322258	2+0-	20	40322449	0+2-	INS	-132	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40324646	2+2-	20	40324606	2+2-	INS	-390	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40330322	2+2-	20	40330331	2+2-	INS	-237	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40335981	2+2-	20	40335992	2+2-	INS	-105	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40350624	2+2-	20	40350584	2+2-	INS	-389	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40361117	2+0-	20	40361138	1+3-	INS	-295	27	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	40387896	2+0-	20	40388031	0+2-	INS	-192	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40401631	2+2-	20	40401645	2+2-	INS	-221	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40404744	2+2-	20	40404706	2+2-	INS	-107	37	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40433542	2+4-	20	40433590	2+4-	INS	-207	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40441452	2+2-	20	40441471	2+2-	INS	-95	29	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40448242	2+2-	20	40448290	2+4-	INS	-120	34	4	COLO-829BL-IL|2:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40451554	2+2-	20	40451525	2+2-	INS	-114	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40458362	2+2-	20	40458395	2+2-	INS	-97	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40476440	2+2-	20	40476438	2+2-	INS	-235	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40479046	2+2-	20	40479038	2+2-	INS	-115	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40483839	3+2-	20	40483904	3+2-	INS	-104	21	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40494189	2+4-	20	40494237	2+4-	INS	-238	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40508575	2+2-	20	40508533	2+2-	INS	-104	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40533291	4+1-	20	40533380	0+3-	INS	-201	41	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	40539011	4+4-	20	40539163	4+4-	INS	-192	21	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40555154	3+3-	20	40555153	3+3-	INS	-282	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40568385	2+0-	20	40569154	2+0-	INV	657	60	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40571830	4+2-	20	40571875	4+2-	INS	-87	26	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40575322	2+3-	20	40575342	2+3-	INS	-100	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40585319	2+0-	20	40585485	0+2-	INS	-163	24	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	40595042	2+1-	20	40595107	0+2-	INS	-227	16	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	40596915	2+2-	20	40596902	2+2-	INS	-257	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40603462	2+2-	20	40603474	2+2-	INS	-218	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40613431	2+2-	20	40613399	2+2-	INS	-111	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40627870	4+1-	20	40627865	1+3-	INS	-220	40	4	COLO-829_v2_74|2:COLO-829-IL|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	40630521	2+2-	20	40630490	2+2-	INS	-120	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40632800	2+2-	20	40632803	2+2-	INS	-108	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40639798	2+0-	20	40639939	3+6-	INS	-92	43	3	COLO-829BL-IL|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	40651585	2+2-	20	40651608	2+2-	INS	-99	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40666096	4+1-	20	40666096	0+3-	INS	-252	40	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	40696524	2+0-	20	40696560	1+3-	INS	-316	32	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	40699558	2+2-	20	40699549	2+2-	INS	-100	32	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40705278	2+0-	20	40705330	3+5-	INS	-177	34	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	40731923	3+3-	20	40731896	3+3-	INS	-115	46	3	COLO-829BL-IL|1:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	40756129	2+2-	20	40756148	2+2-	INS	-108	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40762263	3+0-	20	40762251	0+2-	INS	-345	26	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	40762673	2+2-	20	40762681	2+2-	INS	-89	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40773057	3+0-	20	40773157	1+4-	INS	-202	38	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40792695	3+3-	20	40792743	3+3-	INS	-232	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40805291	2+3-	20	40805415	2+3-	INS	-188	14	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40809738	2+2-	20	40809759	2+2-	INS	-107	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40815292	2+2-	20	40815293	2+2-	INS	-97	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40836120	3+2-	20	40836099	3+2-	INS	-118	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40843127	5+5-	20	40843171	5+5-	INS	-252	48	5	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	40866987	3+3-	20	40867054	1+3-	INS	-207	31	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40906494	2+2-	20	40906503	2+2-	INS	-245	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40923693	3+3-	20	40923782	3+3-	INS	-96	32	3	COLO-829BL-IL|2:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	40931301	3+0-	20	40931354	0+3-	INS	-274	33	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	40945731	4+2-	20	40945794	4+2-	INS	-207	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40945864	2+0-	20	40945875	0+2-	DEL	91	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40952926	2+3-	20	40952876	2+3-	INS	-117	36	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	40959942	2+2-	20	40959937	2+2-	INS	-106	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	40979835	2+0-	20	40979914	1+3-	INS	-193	32	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	41002676	6+2-	20	41002793	6+2-	INS	-254	14	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41004324	2+2-	20	41004284	2+2-	INS	-111	34	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	41008733	3+3-	20	41008747	3+3-	INS	-403	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41020331	2+2-	20	41020365	2+2-	INS	-90	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	41029468	2+2-	20	41029451	2+2-	INS	-87	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41030240	3+1-	20	41030344	0+3-	INS	-161	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	41031339	2+2-	20	41031318	2+2-	INS	-109	34	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	41045972	2+2-	20	41046007	2+2-	INS	-362	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41047617	3+3-	20	41047599	3+3-	INS	-105	44	3	COLO-829BL-IL|1:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	41087776	2+2-	20	41087794	2+2-	INS	-374	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41102762	2+0-	20	41102914	0+2-	INS	-167	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41125536	2+2-	20	41125541	2+2-	INS	-96	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	41127901	3+4-	20	41128025	3+4-	INS	-232	19	3	COLO-829_v2_74|2:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	41158012	6+2-	20	41158066	0+4-	DEL	89	75	4	COLO-829-IL|4	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	41172607	2+2-	20	41172627	2+2-	INS	-116	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41175467	2+2-	20	41175453	2+2-	INS	-105	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	41189985	2+2-	20	41189985	2+2-	INS	-248	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41208292	2+2-	20	41208263	2+2-	INS	-93	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	41213729	3+2-	20	41213710	3+2-	INS	-106	33	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	41218247	2+3-	20	41218334	2+3-	INS	-219	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41219820	3+0-	20	41219890	0+3-	INS	-242	32	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	41229309	2+2-	20	41229338	2+2-	INS	-245	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41234109	2+3-	20	41234126	2+3-	INS	-107	29	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41238309	2+0-	20	41238349	0+2-	INS	-294	26	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	41272556	2+1-	20	41272746	1+3-	INS	-115	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	41276375	2+0-	20	41276371	2+3-	INS	-261	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	41286765	2+2-	20	41286772	2+2-	INS	-96	30	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	41317062	2+2-	20	41317031	2+2-	INS	-102	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41331469	2+2-	20	41331463	2+2-	INS	-248	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41331641	2+2-	20	41331599	2+2-	INS	-104	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41333323	2+2-	20	41333335	2+2-	INS	-94	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	41362283	2+2-	20	41362276	2+2-	INS	-104	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41381933	2+2-	20	41381947	2+2-	INS	-222	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41382881	2+3-	20	41382853	2+3-	INS	-108	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41386390	3+3-	20	41386361	3+3-	INS	-111	49	3	COLO-829BL-IL|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	41399036	2+2-	20	41399049	2+2-	INS	-104	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	41429633	2+3-	20	41429618	2+3-	INS	-97	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41438553	2+2-	20	41438515	2+2-	INS	-254	28	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41440583	3+1-	20	41440608	1+2-	INS	-210	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	41457675	2+0-	20	41459207	1+56-	DEL	1219	42	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	41458026	56+1-	20	41459207	0+53-	DEL	1203	99	53	COLO-829BL-IL|16:COLO-829_v2_74|8:COLO-829-IL|29	0.29	BreakDancerMax-0.0.1r81	|q10|o20
20	41458026	2+0-	20	41459530	1+2-	DEL	1193	38	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	41462634	2+2-	20	41462666	2+2-	INS	-233	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41472648	3+0-	20	41472655	1+4-	INS	-229	27	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	41481371	2+3-	20	41481358	2+3-	INS	-107	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	41510540	4+1-	20	41510527	1+5-	INS	-95	76	5	COLO-829BL-IL|2:COLO-829-IL|3	0.28	BreakDancerMax-0.0.1r81	|q10|o20
20	41525699	2+2-	20	41525645	2+2-	INS	-115	37	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41532907	2+2-	20	41532879	2+2-	INS	-95	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	41577982	2+2-	20	41577999	2+2-	INS	-101	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	41590659	2+3-	20	41590646	2+3-	INS	-104	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41616676	2+2-	20	41616648	2+2-	INS	-104	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41655563	3+2-	20	41655641	3+2-	INS	-232	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41681825	3+0-	20	41681872	0+3-	INS	-252	32	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	41689631	3+2-	20	41689651	3+2-	INS	-106	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	41705313	44+0-	20	41708012	1+48-	DEL	2720	99	41	COLO-829BL-IL|10:COLO-829-IL|31	0.67	BreakDancerMax-0.0.1r81	|q10|o20
20	41731955	3+3-	20	41731974	3+3-	INS	-109	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	41743288	2+2-	20	41743288	2+2-	INS	-100	27	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	41758904	12+48-	20	41758902	39+3-	ITX	6	99	45	COLO-829BL-IL|13:COLO-829_v2_74|9:COLO-829-IL|23	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	41782020	2+2-	20	41781971	2+2-	INS	-405	29	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41820422	3+3-	20	41820495	3+3-	INS	-240	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	41823528	2+1-	20	41823739	0+3-	INS	-132	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41834232	2+1-	20	41834307	0+3-	INS	-255	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41836752	2+3-	20	41836795	2+3-	INS	-100	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41840446	2+2-	20	41840436	2+2-	INS	-97	32	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	41871360	3+3-	20	41871337	3+3-	INS	-373	37	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41882619	2+11-	20	41882672	2+11-	INS	-102	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41905230	2+2-	20	41905232	2+2-	INS	-225	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41906616	3+2-	20	41906673	3+2-	INS	-196	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41914721	19+0-	20	41917195	0+17-	DEL	2525	99	16	COLO-829BL-IL|6:COLO-829-IL|10	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	41925116	2+3-	20	41925100	2+3-	INS	-100	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	41962423	3+2-	20	41962461	3+2-	INS	-104	27	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41963083	2+1-	20	41963150	0+2-	INS	-281	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41973536	2+3-	20	41973580	2+3-	INS	-95	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41974897	2+2-	20	41974885	2+2-	INS	-95	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	41982695	2+2-	20	41982649	2+2-	INS	-259	30	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	41991555	2+2-	20	41991565	2+2-	INS	-256	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42000126	2+2-	20	42000146	2+2-	INS	-90	29	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42005012	2+2-	20	42004987	2+2-	INS	-113	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42008804	2+2-	20	42008763	2+2-	INS	-391	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42012608	2+2-	20	42012620	2+2-	INS	-252	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	42019362	2+3-	20	42019361	2+3-	INS	-118	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42028155	3+1-	20	42028268	0+2-	INS	-165	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42040598	2+2-	20	42040591	2+2-	INS	-111	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42046442	2+2-	20	42046426	2+2-	INS	-93	33	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42060320	3+1-	20	42060450	0+4-	INS	-163	31	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	42060434	3+1-	20	42060450	0+2-	INS	-195	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42073153	3+3-	20	42073174	3+3-	INS	-379	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42074983	3+0-	20	42075141	1+3-	INS	-130	32	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	42085069	2+2-	20	42085044	2+2-	INS	-109	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42088681	2+1-	20	42088802	0+2-	INS	-206	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42109564	36+0-	20	42109864	8+30-	DEL	400	99	29	COLO-829BL-IL|15:COLO-829-IL|14	0.28	BreakDancerMax-0.0.1r81	|q10|o20
20	42109564	7+0-	20	42110177	0+5-	DEL	391	99	5	COLO-829_v2_74|5	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	42114033	2+3-	20	42113996	2+3-	INS	-105	33	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42141842	2+2-	20	42141834	2+2-	INS	-109	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42150421	2+3-	20	42150426	2+3-	INS	-111	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42152769	3+4-	20	42152901	3+4-	INS	-237	18	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42161970	2+2-	20	42161941	2+2-	ITX	-130	45	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42171758	2+3-	20	42171716	2+3-	INS	-110	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42243551	2+0-	20	42243696	0+2-	INS	-179	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42251503	2+3-	20	42251541	2+3-	INS	-365	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42276775	2+2-	20	42276739	2+2-	INS	-106	33	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42281194	5+5-	20	42281325	5+5-	INS	-204	36	5	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42293856	3+3-	20	42293857	3+3-	INS	-388	19	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42299194	2+2-	20	42299144	2+2-	INS	-115	36	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42323557	3+0-	20	42323689	0+3-	INS	-194	32	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42324678	2+3-	20	42324691	2+3-	INS	-115	29	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42331690	2+2-	20	42331706	2+2-	INS	-102	25	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42363852	2+2-	20	42363856	2+2-	INS	-215	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42382275	3+1-	20	42382384	0+2-	INS	-159	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42403561	2+2-	20	42403545	2+2-	INS	-115	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42411389	2+2-	20	42411348	2+2-	INS	-391	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42420153	4+1-	20	42420226	1+3-	INS	-174	41	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42434360	2+2-	20	42434334	2+2-	INS	-113	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	42444982	2+4-	20	42445019	2+4-	INS	-229	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42453111	3+4-	20	42453149	3+4-	INS	-250	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42466813	5+1-	20	42466835	5+14-	DEL	91	80	5	COLO-829BL-IL|1:COLO-829-IL|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42477062	2+2-	20	42477032	2+2-	INS	-100	31	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42477380	3+3-	20	42477454	3+3-	INS	-189	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42479293	4+4-	20	42479393	4+4-	INS	-106	42	4	COLO-829BL-IL|2:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42493643	3+2-	20	42493683	3+2-	INS	-389	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42515070	2+2-	20	42515051	2+2-	INS	-117	29	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42538365	2+2-	20	42538374	2+2-	INS	-253	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42550207	3+4-	20	42550239	3+4-	INS	-255	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42576129	2+2-	20	42576194	0+2-	INS	-257	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42583287	3+1-	20	42583414	0+4-	INS	-184	45	3	COLO-829_v2_74|2:COLO-829-IL|1	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	42597913	2+2-	20	42597872	2+2-	ITX	-129	47	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	42622875	4+3-	20	42622854	4+3-	INS	-298	35	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42623937	2+2-	20	42624004	2+2-	INS	-92	25	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42627360	3+2-	20	42627434	3+2-	INS	-224	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42648495	3+4-	20	42648492	3+4-	INS	-112	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42651347	3+0-	20	42651397	0+3-	INS	-257	33	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42653041	2+2-	20	42652984	2+2-	INS	-407	33	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42663569	2+0-	20	42663704	0+2-	INS	-148	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42683864	3+2-	20	42683936	0+3-	INS	-185	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42715627	2+3-	20	42715667	2+3-	INS	-105	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42723738	2+0-	20	42723869	0+2-	INS	-200	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42737229	2+2-	20	42737192	2+2-	INS	-109	33	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	42753023	4+4-	20	42753115	4+4-	INS	-231	31	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42763384	2+3-	20	42763433	2+3-	INS	-241	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42774352	30+11-	20	42774404	30+11-	INS	-94	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42785622	2+2-	20	42785617	2+2-	INS	-103	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42797065	2+0-	20	42797129	1+3-	INS	-206	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42816166	3+2-	20	42816173	3+2-	INS	-247	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42816385	2+3-	20	42816349	2+3-	INS	-254	26	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42825987	52+60-	20	42826591	52+60-	INS	-113	99	33	COLO-829BL-IL|9:COLO-829_v2_74|10:COLO-829-IL|14	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	42846405	3+1-	20	42846508	0+3-	INS	-197	30	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42849402	2+4-	20	42849421	2+4-	INS	-103	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42850540	2+2-	20	42850506	2+2-	INS	-108	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42870712	2+2-	20	42870677	2+2-	INS	-111	32	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42877143	3+0-	20	42877314	0+2-	INS	-159	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42878044	2+2-	20	42878040	2+2-	INS	-116	27	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42897885	2+1-	20	42898019	0+2-	INS	-170	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42901778	2+2-	20	42901758	2+2-	INS	-99	29	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42905416	2+1-	20	42905491	1+3-	INS	-186	21	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42920958	3+3-	20	42921021	3+3-	INS	-110	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42921343	3+4-	20	42921342	3+4-	INS	-101	42	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42923806	3+1-	20	42923908	1+2-	INS	-171	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42926270	3+4-	20	42926352	3+4-	INS	-112	31	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42936556	3+4-	20	42936564	3+4-	INS	-280	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	42937181	3+1-	20	42937395	0+2-	INS	-121	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42940854	2+2-	20	42940847	2+2-	INS	-104	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42945496	4+1-	20	42945642	0+3-	INS	-162	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42946349	3+3-	20	42946410	3+3-	INS	-379	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42949179	2+3-	20	42949178	2+3-	INS	-109	31	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	42958851	2+0-	20	42958947	0+2-	INS	-221	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42959494	2+2-	20	42959513	2+2-	INS	-98	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	42962486	3+1-	20	42962624	0+2-	INS	-148	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	42993213	7+1-	20	42993338	0+7-	DEL	92	99	7	COLO-829BL-IL|3:COLO-829-IL|4	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	42994064	2+2-	20	42994074	2+2-	INS	-105	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43013536	2+2-	20	43013573	2+2-	INS	-95	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43017867	2+1-	20	43018046	0+2-	INS	-153	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43025392	2+0-	20	43025527	1+6-	INS	-116	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	43025510	2+0-	20	43025527	0+3-	INS	-216	14	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43027789	3+0-	20	43027900	0+4-	INS	-180	26	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	43037267	2+3-	20	43037258	2+3-	INS	-397	21	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	43063893	2+0-	20	43064027	0+2-	INS	-185	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43071920	2+2-	20	43071942	2+2-	INS	-242	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	43075893	2+2-	20	43075866	2+2-	INS	-376	23	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	43083536	2+2-	20	43083546	2+2-	INS	-93	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43097718	3+3-	20	43097804	3+3-	INS	-252	23	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43123171	3+2-	20	43123200	3+2-	INS	-103	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43130830	2+1-	20	43130949	0+3-	INS	-230	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43141138	3+2-	20	43141147	3+2-	INS	-96	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43151740	4+2-	20	43151806	0+2-	INS	-251	45	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	43155942	2+2-	20	43155960	2+2-	INS	-104	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43162652	2+0-	20	43162684	2+4-	INS	-279	37	4	COLO-829_v2_74|4	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	43203798	2+1-	20	43203886	1+2-	INS	-240	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43221780	2+2-	20	43221746	2+2-	INS	-102	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43223933	2+2-	20	43223913	2+2-	INS	-114	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43235226	2+2-	20	43235247	2+2-	INS	-213	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43246664	3+7-	20	43246765	3+7-	INS	-115	19	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43260579	2+0-	20	43260690	2+3-	INS	-230	26	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43280022	2+3-	20	43280060	2+3-	INS	-96	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43317593	2+2-	20	43317605	2+2-	INS	-98	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43325054	2+0-	20	43325166	1+3-	INS	-181	37	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43332749	2+3-	20	43332760	2+3-	INS	-385	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43333845	2+0-	20	43334025	0+2-	INS	-136	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43345818	2+2-	20	43345806	2+2-	INS	-119	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	43363566	2+2-	20	43363560	2+2-	INS	-105	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43371880	3+3-	20	43371978	3+3-	INS	-154	24	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43372242	2+2-	20	43372196	2+2-	INS	-115	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	43403528	2+0-	20	43403625	0+2-	INS	-219	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43413889	4+2-	20	43413876	4+2-	INS	-382	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43417256	2+2-	20	43417260	2+2-	INS	-91	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	43419477	5+2-	20	43419611	5+2-	INS	-205	11	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43419937	4+3-	20	43420000	4+3-	INS	-197	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43423006	4+3-	20	43423036	4+3-	INS	-249	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43424154	2+2-	20	43424124	2+2-	INS	-246	26	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43430337	2+2-	20	43430303	2+2-	INS	-96	32	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	43432331	2+2-	20	43432303	2+2-	INS	-103	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43435127	2+2-	20	43435102	2+2-	INS	-96	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	43441438	2+2-	20	43441424	2+2-	INS	-100	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43441998	2+2-	20	43442045	2+2-	INS	-195	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43461522	2+0-	20	43461566	0+2-	INS	-268	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43466221	2+0-	20	43466349	1+3-	INS	-166	34	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43470888	2+2-	20	43470968	2+2-	INS	-107	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43473504	2+2-	20	43473468	2+2-	INS	-94	33	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43480983	3+3-	20	43480996	3+3-	INS	-102	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43489666	2+3-	20	43489684	2+3-	INS	-92	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43501031	2+4-	20	43501140	2+4-	INS	-96	17	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43516097	3+0-	20	43516091	1+3-	INS	-295	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43530596	2+2-	20	43530643	2+2-	INS	-88	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43534635	9+0-	20	43534747	1+9-	DEL	95	99	8	COLO-829BL-IL|5:COLO-829-IL|3	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	43551551	3+1-	20	43551750	0+2-	INS	-128	37	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43576617	2+2-	20	43576680	2+2-	INS	-107	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43588026	2+2-	20	43588037	2+2-	INS	-100	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	43593610	2+2-	20	43593601	2+2-	INS	-107	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43598204	2+2-	20	43598208	2+2-	INS	-107	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43604235	2+2-	20	43604230	2+2-	INS	-226	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	43609802	2+2-	20	43609821	2+2-	INS	-105	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43610845	2+2-	20	43610864	2+2-	INS	-96	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43613933	3+0-	20	43613943	0+3-	INS	-268	25	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43633150	2+1-	20	43633187	0+2-	INS	-278	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43635629	2+2-	20	43635629	2+2-	INS	-226	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43640326	2+2-	20	43640333	2+2-	INS	-91	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	43641524	2+1-	20	43641749	0+2-	INS	-111	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43645344	2+2-	20	43645292	2+2-	INS	-402	31	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43662735	10+8-	20	43662837	10+8-	INS	-97	84	7	COLO-829BL-IL|3:COLO-829-IL|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	43664079	3+3-	20	43664059	3+3-	INS	-206	39	3	COLO-829_v2_74|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43666665	2+0-	20	43666857	0+2-	INS	-127	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43673904	2+2-	20	43673907	2+2-	INS	-101	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43710599	3+3-	20	43710617	3+3-	INS	-94	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	43715000	2+2-	20	43714986	2+2-	INS	-108	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43738605	2+2-	20	43738579	2+2-	INS	-106	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43747004	3+2-	20	43747096	3+2-	INS	-177	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43749681	4+2-	20	43749709	5+5-	INS	-173	49	6	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	43763794	2+0-	20	43763780	1+3-	INS	-174	31	3	COLO-829_v2_74|1:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	43792869	19+1-	20	43792897	0+15-	DEL	94	99	14	COLO-829BL-IL|6:COLO-829-IL|8	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	43792869	5+1-	20	43793144	5+4-	DEL	106	87	4	COLO-829_v2_74|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	43800968	14+3-	20	43801191	72+75-	INS	-109	99	50	COLO-829BL-IL|17:COLO-829-IL|33	0.56	BreakDancerMax-0.0.1r81	|q10|o20
20	43800968	11+2-	20	43801003	1+11-	DEL	104	99	11	COLO-829BL-IL|2:COLO-829-IL|9	0.22	BreakDancerMax-0.0.1r81	|q10|o20
20	43801749	3+3-	20	43801832	3+3-	INS	-226	24	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43821298	4+3-	20	43821369	4+3-	INS	-97	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	43830698	2+0-	20	43830895	0+2-	INS	-112	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43835735	4+1-	20	43836024	0+52-	DEL	133	90	4	COLO-829_v2_74|4	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	43835914	47+1-	20	43836024	0+48-	DEL	123	99	46	COLO-829BL-IL|15:COLO-829-IL|31	0.79	BreakDancerMax-0.0.1r81	|q10|o20
20	43838164	2+0-	20	43838240	0+2-	INS	-246	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43841157	2+2-	20	43841167	2+2-	INS	-253	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43854954	2+3-	20	43854912	2+3-	INS	-406	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43873447	2+1-	20	43873437	0+2-	INS	-336	23	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	43917916	2+2-	20	43917946	2+2-	INS	-91	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43941891	2+2-	20	43941866	2+2-	INS	-115	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43949892	5+3-	20	43950005	5+3-	INS	-110	19	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	43966572	3+3-	20	43966602	3+3-	INS	-371	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43968811	14+1-	20	43969183	0+13-	DEL	444	99	13	COLO-829BL-IL|4:COLO-829-IL|9	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	43983980	3+1-	20	43984145	2+2-	INS	-156	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	43986733	4+3-	20	43986792	4+3-	INS	-254	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	43989569	3+2-	20	43989596	3+2-	INS	-103	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	43992505	4+3-	20	43992542	4+3-	INS	-191	30	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44004069	347+7-	20	44004043	347+7-	INS	-101	99	6	COLO-829BL-IL|2:COLO-829-IL|4	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44013602	2+3-	20	44013603	2+3-	INS	-372	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44015557	3+4-	20	44015566	0+2-	INS	-302	24	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44057853	8+2-	20	44057837	8+2-	ITX	-130	42	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44085946	2+2-	20	44085932	2+2-	INS	-249	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44110979	2+2-	20	44110984	2+2-	INS	-108	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44128979	3+1-	20	44129032	2+2-	INS	-228	34	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	44138387	3+1-	20	44138436	0+2-	INS	-160	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44143013	2+2-	20	44143023	2+2-	INS	-96	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44147945	2+0-	20	44147926	2+5-	INS	-160	17	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	44150121	2+2-	20	44150137	2+2-	INS	-98	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44170557	2+2-	20	44170538	2+2-	INS	-96	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44204060	2+1-	20	44204077	0+3-	INS	-252	13	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44209651	2+2-	20	44209657	2+2-	INS	-88	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44213522	2+0-	20	44213583	0+2-	INS	-271	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44237920	2+2-	20	44237982	0+2-	INS	-214	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44245704	2+0-	20	44245696	1+3-	INS	-245	30	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	44290072	2+2-	20	44290022	2+2-	INS	-118	36	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	44291610	2+2-	20	44291616	2+2-	INS	-111	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44293030	2+0-	20	44293079	0+2-	INS	-263	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44300986	2+3-	20	44300975	2+3-	INS	-238	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44305359	2+2-	20	44305390	2+2-	INS	-247	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44325280	2+2-	20	44325222	2+2-	INS	-118	41	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	44334926	2+0-	20	44335025	4+3-	INS	-184	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44335190	3+0-	20	44335187	0+3-	INS	-326	24	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44341516	2+0-	20	44341504	1+3-	INS	-189	40	3	COLO-829_v2_74|1:COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	44345936	2+2-	20	44345918	2+2-	INS	-85	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44362559	2+1-	20	44362572	0+3-	INS	-275	20	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	44383009	2+0-	20	44383196	0+2-	INS	-136	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44402133	2+3-	20	44402136	2+3-	INS	-238	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	44412252	2+2-	20	44412273	2+2-	INS	-99	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44430684	2+1-	20	44430715	0+2-	INS	-260	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44441838	2+3-	20	44441833	2+3-	INS	-123	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44458412	2+2-	20	44458417	2+2-	INS	-97	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44465747	4+2-	20	44465755	4+2-	INS	-110	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44474206	3+3-	20	44474248	3+3-	INS	-91	23	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44481086	2+1-	20	44481164	0+2-	INS	-251	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44486863	2+2-	20	44486899	2+2-	INS	-91	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	44520737	2+0-	20	44520923	0+2-	INS	-143	24	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	44526038	2+0-	20	44526124	0+2-	INS	-238	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44529010	2+2-	20	44529024	2+2-	INS	-108	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44532390	2+2-	20	44532430	2+2-	INS	-221	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44537062	2+3-	20	44537089	2+3-	INS	-92	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44537767	2+4-	20	44537793	2+4-	INS	-103	24	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	44557561	2+2-	20	44557529	2+2-	INS	-102	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	44563285	2+2-	20	44563273	2+2-	INS	-88	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44576581	2+3-	20	44576630	2+3-	INS	-109	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44590871	2+2-	20	44590839	2+2-	INS	-102	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	44593934	2+2-	20	44593965	2+2-	INS	-238	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44612908	3+2-	20	44612914	3+2-	INS	-94	30	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44639070	18+1-	20	44639130	39+56-	INS	-112	99	22	COLO-829BL-IL|8:COLO-829-IL|14	0.16	BreakDancerMax-0.0.1r81	|q10|o20
20	44644944	2+0-	20	44645003	0+2-	INS	-258	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44645367	2+0-	20	44645547	1+3-	INS	-135	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44661353	2+2-	20	44661335	2+2-	INS	-368	22	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	44699461	3+3-	20	44699477	3+3-	INS	-180	31	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44703290	3+1-	20	44703434	0+2-	INS	-182	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44704235	2+3-	20	44704286	2+3-	INS	-342	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44707120	2+1-	20	44707238	0+2-	INS	-162	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44709668	2+2-	20	44709678	2+2-	INS	-253	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44740738	3+0-	20	44740821	0+4-	INS	-198	26	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44754563	2+2-	20	44754616	2+2-	INS	-249	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44767077	2+2-	20	44767032	2+2-	INS	-112	35	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44786839	3+3-	20	44786811	3+3-	INS	-86	56	3	COLO-829BL-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44790423	2+2-	20	44790428	2+2-	INS	-225	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44801887	2+1-	20	44802041	0+2-	INS	-140	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44850852	2+1-	20	44850875	76+78-	DEL	98	99	48	COLO-829BL-IL|21:COLO-829_v2_74|2:COLO-829-IL|25	0.54	BreakDancerMax-0.0.1r81	|q10|o20
20	44855105	2+1-	20	44855129	0+2-	INS	-298	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44873958	3+4-	20	44873998	3+4-	INS	-104	37	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44884665	2+3-	20	44884634	2+3-	INS	-100	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44890205	2+3-	20	44890260	2+3-	INS	-94	26	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44893888	4+1-	20	44893870	1+4-	INS	-208	40	5	COLO-829_v2_74|3:COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	44895340	3+1-	20	44895360	0+2-	INS	-230	31	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44902263	2+2-	20	44902286	2+2-	INS	-101	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44912837	2+2-	20	44912836	2+2-	INS	-239	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	44936745	2+3-	20	44936756	2+3-	INS	-99	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	44958575	3+3-	20	44958540	3+3-	INS	-290	42	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44965424	2+1-	20	44965544	0+2-	INS	-183	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44974439	3+3-	20	44974445	3+3-	INS	-112	39	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44978516	2+2-	20	44978496	2+2-	INS	-106	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44980693	3+0-	20	44980682	0+2-	INS	-339	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	44980962	3+3-	20	44981046	3+3-	INS	-186	25	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44983483	3+3-	20	44983489	3+3-	INS	-113	39	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	44989937	2+1-	20	44989918	0+2-	INS	-327	19	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	45010947	2+2-	20	45010936	2+2-	INS	-87	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45012046	2+2-	20	45012061	2+2-	INS	-218	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	45022127	2+3-	20	45022141	2+3-	INS	-236	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45024993	2+0-	20	45025043	0+3-	INS	-240	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45033884	2+2-	20	45033841	2+2-	INS	-111	35	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45039671	2+2-	20	45039684	2+2-	INS	-224	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45044095	2+2-	20	45044093	2+2-	INS	-92	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45066034	2+2-	20	45066011	2+2-	INS	-109	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45070022	2+0-	20	45070009	0+2-	INS	-344	25	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	45094265	3+5-	20	45094436	3+5-	INS	-285	18	3	COLO-829_v2_74|3	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	45107249	2+2-	20	45107250	2+2-	INS	-250	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45117148	2+0-	20	45117309	0+3-	INS	-156	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45125639	2+0-	20	45125691	0+2-	INS	-267	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45125876	2+2-	20	45125863	2+2-	INS	-251	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45142086	3+3-	20	45142119	3+3-	INS	-283	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45152907	2+2-	20	45152946	2+2-	INS	-213	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45168210	2+2-	20	45168235	2+2-	INS	-363	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45177282	2+3-	20	45177336	2+3-	INS	-91	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	45182827	2+3-	20	45182829	2+3-	INS	-107	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45186280	3+3-	20	45186310	3+3-	INS	-238	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45202034	2+3-	20	45202082	2+3-	INS	-112	22	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	45205302	3+1-	20	45205411	0+3-	INS	-154	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45214967	2+2-	20	45214954	2+2-	INS	-105	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45235091	2+3-	20	45235048	2+3-	INS	-119	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45242117	15+2-	20	45242190	15+2-	INS	-225	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45245074	2+2-	20	45245048	2+2-	INS	-375	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45258631	3+2-	20	45258684	3+2-	INS	-192	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	45276449	2+0-	20	45276439	2+4-	INS	-145	46	4	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|1	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	45291909	3+2-	20	45291916	3+2-	INS	-115	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45299145	3+3-	20	45299210	3+3-	INS	-249	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	45319751	2+2-	20	45319773	2+2-	INS	-90	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45331460	3+3-	20	45331517	3+3-	INS	-98	42	3	COLO-829BL-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45357590	2+2-	20	45357562	2+2-	INS	-96	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45393711	2+2-	20	45393661	2+2-	INS	-111	36	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45410141	4+5-	20	45410238	4+5-	INS	-175	36	4	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45412505	2+2-	20	45412515	2+2-	INS	-98	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45442825	3+4-	20	45442807	3+4-	INS	-105	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45452465	11+0-	20	45452765	3+13-	DEL	338	99	11	COLO-829BL-IL|4:COLO-829-IL|7	0.31	BreakDancerMax-0.0.1r81	|q10|o20
20	45480435	2+2-	20	45480478	2+2-	INS	-101	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45501523	2+2-	20	45501500	2+2-	INS	-92	34	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45519575	2+2-	20	45519532	2+2-	INS	-101	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	45559980	2+0-	20	45559982	3+2-	INS	-319	19	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	45583272	2+2-	20	45583308	2+2-	INS	-202	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45595869	2+2-	20	45595850	2+2-	INS	-247	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45660093	3+0-	20	45660643	2+2-	INV	494	51	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45666690	2+2-	20	45666646	2+2-	INS	-109	35	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45667539	2+2-	20	45667544	2+2-	INS	-107	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	45669433	2+3-	20	45669385	2+3-	INS	-397	29	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45707923	2+2-	20	45707891	2+2-	INS	-99	36	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	45712198	6+2-	20	45712260	6+2-	INS	-241	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45728186	5+0-	20	45728241	19+16-	ITX	-161	99	11	COLO-829BL-IL|2:COLO-829-IL|9	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	45728424	8+0-	20	45728491	0+10-	INS	-167	73	8	COLO-829_v2_74|8	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	45756105	2+2-	20	45756078	2+2-	INS	-250	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45756922	2+3-	20	45756978	2+3-	INS	-104	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45778675	2+4-	20	45778765	2+4-	INS	-207	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45784233	3+2-	20	45784292	3+2-	INS	-189	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45792318	2+2-	20	45792303	2+2-	INS	-123	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45794134	2+0-	20	45794205	0+2-	INS	-231	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45804847	2+0-	20	45805009	0+5-	INS	-158	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45813272	3+1-	20	45813481	0+2-	INS	-117	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	45828353	4+0-	20	45828400	0+4-	INS	-286	61	4	COLO-829_v2_74|4	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	45828815	3+1-	20	45828823	0+2-	INS	-249	35	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	45833058	2+0-	20	45833105	0+2-	INS	-264	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45838224	2+1-	20	45838404	1+2-	INS	-134	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45860385	2+2-	20	45860377	2+2-	INS	-109	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45901021	8+0-	20	45952387	8+0-	INV	51275	99	8	COLO-829BL-IL|4:COLO-829-IL|4	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	45905017	4+14-	20	45974700	8+1-	INV	69616	99	4	COLO-829BL-IL|2:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	45905017	0+14-	20	45974881	0+29-	INV	69840	99	14	COLO-829BL-IL|5:COLO-829-IL|9	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	45907428	2+3-	20	45972637	1+2-	INV	65127	61	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45907428	2+1-	20	45972435	8+2-	INV	64897	47	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45910222	2+2-	20	45910276	2+2-	INS	-232	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45914572	2+2-	20	45914573	2+2-	INS	-251	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45956831	6+0-	20	45956859	495+414-	DEL	96	99	163	COLO-829BL-IL|67:COLO-829_v2_74|1:COLO-829-IL|95	0.39	BreakDancerMax-0.0.1r81	|q10|o20
20	45957655	233+146-	20	45957657	80+93-	DEL	293	99	42	COLO-829BL-IL|16:COLO-829_v2_74|5:COLO-829-IL|21	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45992552	2+2-	20	45992552	2+2-	INS	-259	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45997633	3+0-	20	45997679	1+3-	INS	-228	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46007028	2+0-	20	46007076	0+2-	INS	-261	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46013477	9+9-	20	46013562	9+9-	INS	-103	79	6	COLO-829-IL|6	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46042829	2+2-	20	46042786	2+2-	INS	-392	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46052568	2+3-	20	46052578	2+3-	INS	-243	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46053362	2+2-	20	46053380	2+2-	INS	-107	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46061064	2+0-	20	46061111	1+2-	INS	-276	22	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46061514	2+3-	20	46061517	2+3-	INS	-387	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46066036	4+5-	20	46066143	4+5-	INS	-277	29	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46073157	43+8-	20	46073140	3+37-	INS	-146	99	22	COLO-829_v2_74|18:COLO-829-IL|4	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	46073413	2+1-	20	46073455	0+2-	INS	-118	10	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46125875	3+1-	20	46126000	0+2-	INS	-162	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46132597	2+2-	20	46132633	2+2-	INS	-119	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46134982	2+2-	20	46135006	2+2-	INS	-97	28	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46144035	2+2-	20	46144040	2+2-	INS	-234	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46168263	2+0-	20	46168387	0+2-	INS	-193	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	45897800	8+7-	20	46189666	0+8-	DEL	291854	99	8	COLO-829BL-IL|2:COLO-829-IL|6	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	45897800	0+7-	20	46189402	8+1-	ITX	291458	99	7	COLO-829BL-IL|5:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	46207305	2+0-	20	46207470	0+2-	INS	-159	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46208032	2+2-	20	46208087	0+2-	INS	-229	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46214467	3+3-	20	46214458	3+3-	INS	-105	44	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46224979	3+2-	20	46224973	3+2-	INS	-115	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46226042	2+1-	20	46226230	1+3-	INS	-144	34	3	COLO-829_v2_74|2:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	46236266	2+2-	20	46236213	2+2-	INS	-114	37	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46265395	2+0-	20	46265481	1+3-	INS	-226	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46087219	0+2-	20	46382699	0+2-	INV	295410	51	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46306392	3+1-	20	46306411	1+3-	INS	-205	41	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46307354	4+3-	20	46307399	4+3-	INS	-109	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46335593	2+0-	20	46335673	11+3-	INS	-250	14	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	46337022	2+2-	20	46337001	2+2-	INS	-122	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46338237	2+3-	20	46338218	2+3-	INS	-254	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46349266	2+0-	20	46349348	1+3-	INS	-189	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46358823	2+3-	20	46358832	2+3-	INS	-223	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46369310	2+2-	20	46369283	2+2-	INS	-102	35	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46371747	2+2-	20	46371704	2+2-	INS	-105	39	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46398252	2+0-	20	46398280	0+2-	INS	-292	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46409937	2+2-	20	46409919	2+2-	INS	-105	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46422639	2+1-	20	46422635	0+2-	INS	-180	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46433737	2+2-	20	46433699	2+2-	INS	-387	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46440228	3+0-	20	46440279	1+4-	INS	-206	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46445192	4+3-	20	46445213	4+3-	INS	-101	40	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46453230	10+11-	20	46453420	10+11-	INS	-92	72	7	COLO-829BL-IL|3:COLO-829-IL|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46453490	3+4-	20	46453483	0+2-	INS	-246	8	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46469114	3+3-	20	46469085	3+3-	INS	-100	56	3	COLO-829BL-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	45911398	13+10-	20	46521294	11+1-	ITX	609762	99	10	COLO-829BL-IL|1:COLO-829-IL|9	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	45911398	13+0-	20	46521565	0+13-	DEL	610154	99	13	COLO-829BL-IL|3:COLO-829-IL|10	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	45957655	195+138-	20	46564756	1717+1634-	ITX	132	99	682	COLO-829BL-IL|256:COLO-829_v2_74|94:COLO-829-IL|332	0.25	BreakDancerMax-0.0.1r81	|q10|o20
20	45958267	52+35-	20	46564756	99+76-	INV	607489	99	80	COLO-829BL-IL|32:COLO-829_v2_74|9:COLO-829-IL|39	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	46187655	3+0-	20	46564756	49+44-	DEL	377478	41	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	46188419	3+5-	20	46564756	49+41-	ITX	376761	82	5	COLO-829_v2_74|4:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	45964972	22+15-	20	46557615	2+15-	INV	592600	99	15	COLO-829BL-IL|10:COLO-829-IL|5	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	45964972	22+0-	20	46557360	23+0-	INV	592319	99	22	COLO-829BL-IL|7:COLO-829-IL|15	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	45974828	4+1-	20	46547536	4+15-	INV	572633	99	4	COLO-829BL-IL|2:COLO-829-IL|2	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	45975070	0+15-	20	46547536	0+15-	INV	572390	99	15	COLO-829BL-IL|3:COLO-829-IL|12	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	46475338	2+0-	20	46475450	0+2-	INS	-221	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46480315	2+3-	20	46480298	2+3-	INS	-119	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46482241	2+4-	20	46482291	2+4-	INS	-107	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46488319	3+0-	20	46488377	0+2-	INS	-253	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46493443	22+8-	20	46493571	6+3-	DEL	90	54	3	COLO-829BL-IL|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46493443	19+8-	20	46493424	9+0-	ITX	-162	99	6	COLO-829BL-IL|2:COLO-829-IL|4	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	46493443	19+2-	20	46493793	3+28-	DEL	340	99	19	COLO-829BL-IL|6:COLO-829_v2_74|6:COLO-829-IL|7	0.17	BreakDancerMax-0.0.1r81	|q10|o20
20	46493668	6+0-	20	46493793	1+9-	DEL	135	99	6	COLO-829BL-IL|3:COLO-829-IL|3	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	46493539	3+0-	20	46493793	1+3-	DEL	101	64	3	COLO-829_v2_74|3	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	46495919	3+0-	20	46496065	1+4-	INS	-129	37	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46497717	2+2-	20	46497722	2+2-	INS	-105	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46500383	2+0-	20	46500602	0+2-	INS	-109	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46501180	2+0-	20	46501330	0+3-	INS	-184	21	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46507446	3+3-	20	46507468	3+3-	INS	-105	40	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46511799	15+3-	20	46511966	15+3-	INS	-296	10	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46519640	2+2-	20	46519599	2+2-	INS	-248	27	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46548688	3+2-	20	46548654	3+2-	INS	-255	25	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46276816	0+13-	20	46647953	2+13-	INV	371140	99	13	COLO-829BL-IL|4:COLO-829-IL|9	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	46593788	2+2-	20	46593768	2+2-	INS	-111	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46616540	3+3-	20	46616570	3+3-	INS	-284	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46622056	3+2-	20	46622077	3+2-	INS	-254	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46624212	2+1-	20	46624208	0+3-	INS	-333	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46663063	2+2-	20	46663029	2+2-	INS	-383	25	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46672916	3+3-	20	46672964	3+3-	INS	-93	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46691817	16+6-	20	46691831	16+6-	INS	-91	40	3	COLO-829BL-IL|2:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	46724670	2+2-	20	46724706	2+2-	INS	-246	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46739945	3+2-	20	46739930	3+2-	INS	-380	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46761101	2+2-	20	46761076	2+2-	INS	-374	23	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46796446	2+2-	20	46796461	2+2-	INS	-230	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46801385	2+2-	20	46801393	2+2-	INS	-98	30	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46827838	4+0-	20	46827949	0+4-	INS	-189	39	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46843454	2+0-	20	46843580	0+2-	INS	-194	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46846081	2+3-	20	46846072	2+3-	INS	-101	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	46847446	2+2-	20	46847434	2+2-	INS	-91	28	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46858715	2+0-	20	46858941	1+2-	INS	-106	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46867418	2+2-	20	46867418	2+2-	INS	-245	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46872728	2+0-	20	46872875	0+2-	INS	-170	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46874889	2+0-	20	46874935	0+3-	INS	-238	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46880644	2+2-	20	46880614	2+2-	INS	-119	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46880843	2+2-	20	46880864	2+2-	INS	-102	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46882793	2+2-	20	46882820	2+2-	INS	-212	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46889290	3+3-	20	46889296	3+3-	INS	-113	41	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46889628	4+3-	20	46889681	4+3-	INS	-175	26	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46901904	3+2-	20	46901980	3+2-	INS	-96	24	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46902362	3+1-	20	46902428	1+3-	INS	-173	44	4	COLO-829_v2_74|2:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46906139	2+0-	20	46906134	0+3-	INS	-295	15	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46907191	2+0-	20	46907280	1+3-	INS	-227	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46927374	2+2-	20	46927327	2+2-	INS	-105	40	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46946678	2+2-	20	46946654	2+2-	INS	-373	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	46947165	17+9-	20	46947212	17+9-	INS	-94	22	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	46974903	2+2-	20	46974929	2+2-	INS	-99	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46989413	2+0-	20	46989487	0+2-	INS	-231	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	46994017	3+1-	20	46994082	2+3-	INS	-228	36	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	47004201	2+2-	20	47004204	2+2-	INS	-116	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47017493	2+4-	20	47017573	2+4-	INS	-188	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47019254	3+2-	20	47019257	3+2-	INS	-373	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47039388	2+2-	20	47039330	2+2-	INS	-408	34	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	47041728	3+1-	20	47041717	0+2-	INS	-319	27	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	47052297	2+2-	20	47052266	2+2-	INS	-380	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47063303	2+0-	20	47063421	0+2-	INS	-208	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47064889	4+2-	20	47064968	4+2-	INS	-95	24	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47079635	2+2-	20	47079623	2+2-	INS	-117	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	47101512	2+2-	20	47101470	2+2-	INS	-106	38	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47102029	2+0-	20	47102018	3+3-	INS	-212	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	47102211	2+0-	20	47102256	0+2-	INS	-176	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47112870	2+2-	20	47112912	2+2-	INS	-240	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47119212	2+0-	20	47119338	0+2-	INS	-184	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47119781	2+2-	20	47119743	2+2-	INS	-107	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47142144	3+3-	20	47142162	3+3-	INS	-93	39	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47156644	3+2-	20	47156658	3+2-	INS	-100	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47157172	2+0-	20	47157223	2+3-	INS	-200	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	47163655	2+3-	20	47163709	2+3-	INS	-203	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47185927	2+5-	20	47186072	2+5-	INS	-237	13	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	47209226	2+2-	20	47209192	2+2-	INS	-91	36	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	47210206	2+2-	20	47210193	2+2-	INS	-237	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47223605	2+2-	20	47223688	0+4-	INS	-207	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47229465	2+2-	20	47229412	2+2-	INS	-402	31	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47233571	2+0-	20	47233589	0+2-	INS	-291	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47250065	2+0-	20	47250206	2+2-	INS	-149	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47265857	2+3-	20	47265814	2+3-	INS	-112	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47297053	3+1-	20	47297105	1+3-	INS	-185	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	47326141	2+3-	20	47326148	2+3-	INS	-104	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47330283	2+0-	20	47330278	1+3-	INS	-321	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47330671	2+3-	20	47330699	2+3-	INS	-236	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	47332594	2+2-	20	47332546	2+2-	ITX	-126	50	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	47338150	3+0-	20	47338181	3+3-	INS	-266	18	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47395608	2+2-	20	47395561	2+2-	INS	-117	40	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47404982	3+0-	20	47405038	0+2-	INS	-266	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47424570	5+0-	20	47424632	1+6-	INS	-191	52	6	COLO-829_v2_74|5:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	47425095	2+2-	20	47425100	2+2-	INS	-94	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47471398	2+2-	20	47471356	2+2-	INS	-99	38	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	47473734	2+2-	20	47473766	2+2-	INS	-247	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47486166	2+3-	20	47486149	2+3-	INS	-369	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47486664	2+4-	20	47486742	2+4-	INS	-91	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	47506216	3+1-	20	47506330	0+2-	INS	-200	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47546634	9+1-	20	47547486	2+14-	DEL	965	99	9	COLO-829BL-IL|3:COLO-829-IL|6	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	47547438	3+0-	20	47547486	0+3-	INS	-130	10	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	47556010	2+2-	20	47555984	2+2-	INS	-102	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47573306	2+2-	20	47573316	2+2-	INS	-99	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47582809	2+2-	20	47582965	1+3-	INS	-128	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47584491	2+2-	20	47584495	2+2-	INS	-91	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47600322	2+2-	20	47600298	2+2-	INS	-100	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47605203	2+1-	20	47605216	1+3-	INS	-99	42	3	COLO-829BL-IL|2:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	47619316	2+2-	20	47619313	2+2-	INS	-231	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47631321	2+2-	20	47631287	2+2-	INS	-383	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47644156	2+2-	20	47644133	2+2-	INS	-95	34	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	47667360	3+0-	20	47667551	8+6-	DEL	166	63	3	COLO-829-IL|3	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	47667561	15+20-	20	47667551	6+1-	ITX	-145	99	13	COLO-829BL-IL|3:COLO-829-IL|10	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	47680503	2+0-	20	47680690	0+3-	INS	-136	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47685025	3+1-	20	47685054	0+2-	INS	-228	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	47692663	2+2-	20	47692679	2+2-	INS	-106	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47708238	2+0-	20	47708295	0+2-	INS	-275	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47719645	3+1-	20	47719636	0+2-	INS	-176	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	47725692	2+2-	20	47725659	2+2-	INS	-245	25	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47734910	2+1-	20	47734990	0+3-	INS	-216	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47759743	2+2-	20	47759714	2+2-	INS	-91	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47771572	3+2-	20	47771680	0+3-	INS	-213	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47793618	3+2-	20	47793643	3+2-	INS	-114	24	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47813268	2+2-	20	47813241	2+2-	INS	-94	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	47842830	2+2-	20	47842886	2+2-	INS	-195	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47893166	2+2-	20	47893202	2+2-	INS	-238	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47906989	3+4-	20	47907044	3+4-	INS	-91	26	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47924295	2+6-	20	47924270	2+6-	INS	-415	23	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	47935498	2+3-	20	47935569	2+3-	INS	-98	25	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	47945026	3+0-	20	47945063	1+3-	INS	-282	35	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47968313	2+1-	20	47968350	0+3-	INS	-223	14	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	47977185	18+1-	20	47977220	0+19-	DEL	95	99	17	COLO-829BL-IL|6:COLO-829-IL|11	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	47995476	4+1-	20	47995507	1+2-	INS	-215	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48011420	2+0-	20	48011438	0+4-	INS	-257	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48013415	1+11-	20	48013397	7+1-	ITX	-83	99	6	COLO-829BL-IL|5:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	48021983	3+3-	20	48022019	3+3-	INS	-110	35	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48036764	2+2-	20	48036728	2+2-	INS	-114	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48041385	2+0-	20	48042350	3+1-	INV	873	52	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	48079101	2+2-	20	48079089	2+2-	INS	-233	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	48084618	2+0-	20	48084811	0+2-	INS	-135	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48111155	2+3-	20	48111130	2+3-	INS	-241	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48123065	2+4-	20	48123086	2+4-	INS	-215	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48159226	3+2-	20	48159189	3+2-	INS	-110	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48178443	2+2-	20	48178398	2+2-	INS	-395	28	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	48184024	5+4-	20	48184067	5+4-	INS	-200	37	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48186984	2+2-	20	48186963	2+2-	INS	-96	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	48192813	3+1-	20	48192842	1+2-	INS	-206	33	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	48193208	2+2-	20	48193164	2+2-	INS	-393	28	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48206219	21+0-	20	48206498	1+18-	DEL	322	99	16	COLO-829BL-IL|7:COLO-829-IL|9	0.28	BreakDancerMax-0.0.1r81	|q10|o20
20	48206219	5+0-	20	48206661	11+2-	DEL	311	42	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	48224553	3+4-	20	48224590	3+4-	INS	-121	23	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48251802	2+2-	20	48251782	2+2-	INS	-102	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	48257189	2+0-	20	48257294	1+4-	INS	-159	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48258563	3+2-	20	48258606	3+2-	INS	-235	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48293723	2+2-	20	48293702	2+2-	INS	-105	30	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	48308107	55+46-	20	48308676	55+46-	INS	-138	99	44	COLO-829BL-IL|7:COLO-829_v2_74|17:COLO-829-IL|20	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	48340095	2+2-	20	48340045	2+2-	INS	-108	36	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	48351086	91+1-	20	48351340	1+8-	DEL	103	99	7	COLO-829_v2_74|7	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	48351086	83+0-	20	48351128	0+83-	DEL	106	99	81	COLO-829BL-IL|25:COLO-829-IL|56	0.49	BreakDancerMax-0.0.1r81	|q10|o20
20	48351086	2+0-	20	48351498	0+2-	DEL	107	42	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48355649	3+3-	20	48355647	3+3-	INS	-279	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48374268	2+1-	20	48374360	0+3-	INS	-153	11	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48398888	3+3-	20	48398907	3+3-	INS	-102	29	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48399794	2+2-	20	48399774	2+2-	INS	-238	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	48409476	3+1-	20	48409527	1+3-	INS	-183	47	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	48416920	2+2-	20	48416954	2+2-	INS	-225	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48451677	2+3-	20	48451648	2+3-	INS	-407	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48466909	2+2-	20	48466932	2+2-	INS	-249	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48467745	2+1-	20	48467946	0+2-	INS	-128	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48484763	2+2-	20	48484798	2+2-	INS	-234	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48532198	2+3-	20	48532200	2+3-	INS	-90	30	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	48538571	3+3-	20	48538542	3+3-	INS	-381	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48552358	3+3-	20	48552399	3+3-	INS	-93	36	3	COLO-829BL-IL|2:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	48561589	3+3-	20	48561604	0+2-	INS	-228	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48563853	2+2-	20	48563847	2+2-	INS	-221	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48565927	2+2-	20	48565894	2+2-	INS	-100	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48570456	3+1-	20	48570567	0+3-	INS	-156	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	48582962	2+6-	20	48583055	2+6-	INS	-374	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48584153	2+2-	20	48584143	2+2-	INS	-224	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48623252	2+2-	20	48623277	2+2-	INS	-93	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	48629596	2+2-	20	48629624	2+2-	INS	-252	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	48639993	2+3-	20	48640027	2+3-	INS	-98	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	48648456	2+0-	20	48648482	1+2-	INS	-246	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48664184	3+2-	20	48664189	3+2-	INS	-97	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48678596	2+2-	20	48678573	2+2-	INS	-92	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48681893	2+0-	20	48681960	0+2-	INS	-253	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48705191	2+2-	20	48705208	2+2-	INS	-232	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48708804	3+1-	20	48708820	0+3-	INS	-320	46	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	48716084	37+24-	20	48716237	37+24-	INS	-93	99	14	COLO-829BL-IL|4:COLO-829-IL|10	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	48733894	5+0-	20	48734121	0+2-	INS	-105	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48784679	2+2-	20	48784676	2+2-	INS	-102	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48794972	3+1-	20	48795044	1+2-	INS	-211	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48802615	2+2-	20	48802606	2+2-	INS	-104	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48808560	2+0-	20	48808732	1+3-	INS	-143	41	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48825774	3+0-	20	48825919	1+3-	DEL	141	61	3	COLO-829-IL|3	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	48827577	2+0-	20	48827614	0+2-	INS	-299	27	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48843465	3+3-	20	48843529	3+3-	INS	-97	35	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48853221	2+1-	20	48853432	1+2-	INS	-137	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48855936	4+2-	20	48856009	4+2-	INS	-101	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48856079	2+0-	20	48856087	0+2-	INS	-180	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48866226	0+21-	20	48866417	35+10-	ITX	129	99	23	COLO-829BL-IL|9:COLO-829_v2_74|3:COLO-829-IL|11	0.17	BreakDancerMax-0.0.1r81	|q10|o20
20	48866412	2+4-	20	48866417	11+6-	ITX	-310	99	4	COLO-829_v2_74|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	48868097	2+2-	20	48868114	2+2-	INS	-96	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48873136	2+4-	20	48873115	2+4-	INS	-114	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48889098	2+2-	20	48889098	2+2-	INS	-379	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48903640	6+1-	20	48903645	9+14-	INS	-152	99	15	COLO-829BL-IL|5:COLO-829_v2_74|7:COLO-829-IL|3	0.16	BreakDancerMax-0.0.1r81	|q10|o20
20	48918834	3+3-	20	48918878	3+3-	INS	-194	29	3	COLO-829_v2_74|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48923429	2+0-	20	48923511	0+2-	INS	-230	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48933972	2+2-	20	48933946	2+2-	INS	-376	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48937217	4+4-	20	48937290	4+4-	INS	-91	33	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48961454	2+0-	20	48961451	1+3-	INS	-102	49	3	COLO-829BL-IL|2:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	48963672	2+2-	20	48963677	2+2-	INS	-92	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	48992516	3+2-	20	48992511	3+2-	INS	-355	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	48995888	2+0-	20	48995876	1+2-	INS	-217	26	2	COLO-829_v2_74|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	48999221	2+2-	20	48999233	2+2-	INS	-217	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49022994	2+2-	20	49022997	2+2-	INS	-95	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49031890	2+3-	20	49031927	2+3-	INS	-97	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49051449	2+2-	20	49051429	2+2-	INS	-110	33	2	COLO-829BL-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	49056555	150+153-	20	49056526	150+153-	INS	-98	99	150	COLO-829BL-IL|56:COLO-829-IL|94	0.23	BreakDancerMax-0.0.1r81	|q10|o20
20	49071699	3+4-	20	49071749	3+4-	INS	-294	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49082438	4+1-	20	49082549	0+2-	INS	-169	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49102317	2+2-	20	49102318	2+2-	INS	-109	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49106028	2+2-	20	49106027	2+2-	INS	-234	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49110945	7+3-	20	49111027	7+3-	INS	-101	20	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49115180	2+2-	20	49115193	2+2-	INS	-89	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49154995	3+2-	20	49154950	3+2-	INS	-112	35	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49163570	5+4-	20	49163644	5+4-	INS	-99	40	3	COLO-829BL-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49207091	2+0-	20	49207269	0+2-	INS	-141	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49218389	2+2-	20	49218362	2+2-	INS	-375	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49223991	2+2-	20	49223987	2+2-	INS	-91	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	49243529	3+2-	20	49243583	3+2-	INS	-105	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49263118	3+1-	20	49263177	0+2-	INS	-244	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49282315	6+2-	20	49282298	6+2-	INS	-233	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	49289841	3+2-	20	49289878	3+2-	INS	-95	27	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49290451	2+3-	20	49290455	2+3-	INS	-102	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49298134	2+0-	20	49298303	0+2-	INS	-171	30	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49300624	2+4-	20	49300689	2+4-	INS	-92	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	49322241	2+1-	20	49322432	3+2-	INS	-131	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49322556	3+0-	20	49322576	1+2-	INS	-259	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49337765	2+0-	20	49337790	0+2-	INS	-271	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49338787	3+0-	20	49338865	1+3-	INS	-212	25	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	49340831	3+2-	20	49340842	3+2-	INS	-99	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49353911	2+2-	20	49353894	2+2-	INS	-113	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	49359137	2+2-	20	49359120	2+2-	INS	-102	33	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49360274	2+2-	20	49360259	2+2-	INS	-103	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49372699	2+0-	20	49372815	1+2-	INS	-196	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49375911	2+0-	20	49376033	0+2-	INS	-195	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49379988	2+2-	20	49379985	2+2-	INS	-114	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49382947	3+0-	20	49383000	1+4-	INS	-256	25	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49390288	2+2-	20	49390289	2+2-	INS	-252	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49403457	2+2-	20	49403450	2+2-	INS	-107	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	49407942	13+12-	20	49407916	13+12-	INS	-119	99	8	COLO-829BL-IL|3:COLO-829-IL|5	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	49407986	2+1-	20	49408095	0+2-	DEL	94	39	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49410159	2+2-	20	49410108	2+2-	INS	-401	30	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	49415589	2+4-	20	49415680	2+4-	INS	-225	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49417560	2+2-	20	49417557	2+2-	INS	-118	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49421577	2+2-	20	49421551	2+2-	INS	-376	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49424563	2+2-	20	49424557	2+2-	INS	-110	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49447317	2+0-	20	49447385	1+3-	INS	-191	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	49457806	2+4-	20	49457804	2+4-	INS	-94	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49465621	2+0-	20	49465712	1+3-	INS	-182	32	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	49475435	3+3-	20	49475428	3+3-	INS	-280	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49480899	2+0-	20	49480978	0+2-	INS	-250	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49484596	3+0-	20	49484598	2+4-	INS	-222	41	4	COLO-829_v2_74|3:COLO-829-IL|1	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	49484818	2+3-	20	49484863	2+3-	INS	-216	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49487129	2+2-	20	49487152	2+2-	INS	-103	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49488970	2+3-	20	49489034	2+3-	INS	-91	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49490246	3+8-	20	49490290	3+8-	INS	-98	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49492937	2+2-	20	49492942	2+2-	INS	-102	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	49511599	2+2-	20	49511604	2+2-	INS	-94	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49517706	2+3-	20	49517788	2+3-	INS	-89	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	49524793	3+3-	20	49524842	3+3-	INS	-93	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49528579	2+2-	20	49528593	2+2-	INS	-254	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49535378	4+4-	20	49535436	4+4-	INS	-222	40	4	COLO-829BL-IL|2:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49579558	2+3-	20	49579538	2+3-	INS	-104	29	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	49593150	2+0-	20	49593207	2+4-	INS	-217	37	4	COLO-829_v2_74|3:COLO-829-IL|1	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	49594954	2+2-	20	49594929	2+2-	INS	-242	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49605101	2+2-	20	49605102	2+2-	INS	-250	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49611798	3+3-	20	49611763	3+3-	INS	-204	42	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49649312	2+2-	20	49649265	2+2-	INS	-111	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49661081	2+0-	20	49661112	2+3-	INS	-303	23	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	49689432	2+0-	20	49689541	1+3-	INS	-169	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	49727425	2+3-	20	49727515	2+3-	INS	-187	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49740765	5+4-	20	49740751	0+2-	INS	-230	37	5	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	49748139	2+0-	20	49748143	0+2-	INS	-308	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49761341	2+2-	20	49761347	2+2-	INS	-102	30	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49772046	2+2-	20	49772014	2+2-	INS	-382	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49790548	6+7-	20	49790541	6+7-	INS	-93	94	6	COLO-829BL-IL|2:COLO-829-IL|4	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	49796234	2+2-	20	49796238	2+2-	INS	-222	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49799813	4+2-	20	49799854	4+2-	INS	-114	23	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49802196	2+4-	20	49802205	2+4-	INS	-95	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49809095	2+0-	20	49809240	0+2-	INS	-194	30	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49828236	3+2-	20	49828227	3+2-	INS	-383	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49894665	3+3-	20	49894715	3+3-	INS	-219	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49896271	2+2-	20	49896233	2+2-	INS	-111	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49898501	2+2-	20	49898467	2+2-	INS	-100	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	49942272	4+2-	20	49942336	4+2-	INS	-206	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49968775	2+1-	20	49968841	0+2-	INS	-237	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	49969858	2+3-	20	49969838	2+3-	ITX	-131	43	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	49970924	2+0-	20	49970965	0+2-	INS	-286	23	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	49975594	22+21-	20	49975632	22+21-	ITX	-141	99	12	COLO-829BL-IL|6:COLO-829-IL|6	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	49982590	2+3-	20	49982570	2+3-	INS	-109	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50001560	6+2-	20	50001635	1+3-	INS	-245	30	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	50002837	2+1-	20	50002829	0+2-	INS	-331	23	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	50004431	2+2-	20	50004452	2+2-	INS	-92	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50025853	3+2-	20	50025825	3+2-	INS	-109	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50029413	2+2-	20	50029392	2+2-	INS	-227	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50043203	3+4-	20	50043251	3+4-	INS	-210	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50056889	2+2-	20	50056878	2+2-	INS	-105	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50063052	2+2-	20	50063076	2+2-	INS	-238	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50064661	2+2-	20	50064621	2+2-	INS	-102	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	50071573	2+3-	20	50071580	2+3-	INS	-110	26	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50072553	2+2-	20	50072566	2+2-	INS	-107	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50103613	3+3-	20	50103777	0+2-	INS	-202	24	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50148408	2+2-	20	50148395	2+2-	INS	-95	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50199695	2+2-	20	50199677	2+2-	INS	-230	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50203770	2+0-	20	50203816	1+3-	INS	-205	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	50207264	4+5-	20	50207371	4+5-	INS	-169	33	4	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50246925	4+1-	20	50246961	1+3-	INS	-174	41	4	COLO-829BL-IL|2:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	50261192	2+2-	20	50261178	2+2-	INS	-233	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50265609	2+1-	20	50265601	2+4-	INS	-227	22	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	50277894	5+3-	20	50278006	5+3-	INS	-109	23	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	50281082	2+2-	20	50281091	2+2-	INS	-222	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50284387	2+2-	20	50284369	2+2-	INS	-98	33	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50320073	2+2-	20	50320028	2+2-	INS	-112	35	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50321905	3+0-	20	50322028	1+2-	INS	-203	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50323581	3+2-	20	50323618	3+2-	INS	-236	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50328318	2+0-	20	50328467	1+3-	INS	-228	28	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50330872	2+3-	20	50330935	2+3-	INS	-97	21	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50340072	2+2-	20	50340069	2+2-	INS	-104	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50351903	2+0-	20	50351945	0+3-	INS	-291	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50353944	2+2-	20	50353989	2+2-	INS	-338	15	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50360579	2+3-	20	50360633	2+3-	INS	-200	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50363726	3+3-	20	50363730	3+3-	INS	-119	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50364892	2+5-	20	50364866	2+5-	INS	-92	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50378868	2+2-	20	50378838	2+2-	INS	-92	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50382894	2+2-	20	50382845	2+2-	INS	-110	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50395598	2+2-	20	50395608	2+2-	INS	-101	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50416063	2+0-	20	50416132	0+2-	INS	-266	27	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50437228	2+2-	20	50437238	2+2-	INS	-109	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50443624	2+2-	20	50443589	2+2-	INS	-92	32	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	50486330	3+3-	20	50486342	3+3-	INS	-90	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50487238	4+3-	20	50487216	4+3-	INS	-109	47	3	COLO-829BL-IL|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	50537719	2+2-	20	50537742	2+2-	INS	-102	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50538453	4+2-	20	50538528	4+2-	INS	-196	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50551816	2+2-	20	50551808	2+2-	INS	-223	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50556390	2+3-	20	50556372	2+3-	INS	-98	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50560754	2+3-	20	50560747	2+3-	INS	-245	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50564723	2+0-	20	50564810	0+2-	INS	-236	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50566254	3+2-	20	50566263	0+2-	INS	-164	26	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50570440	2+2-	20	50570433	2+2-	INS	-92	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50578612	2+2-	20	50578646	2+2-	INS	-96	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50584740	3+1-	20	50584880	1+2-	INS	-115	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50615846	2+0-	20	50615921	0+2-	INS	-240	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50635611	2+3-	20	50635577	2+3-	INS	-101	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50640208	2+2-	20	50640246	2+2-	INS	-199	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50640476	4+4-	20	50640606	4+4-	INS	-199	29	4	COLO-829_v2_74|2:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50647349	3+0-	20	50647398	1+4-	INS	-252	33	4	COLO-829_v2_74|4	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	50651689	2+2-	20	50651642	2+2-	INS	-101	40	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50656240	2+3-	20	50656195	2+3-	INS	-114	39	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50660571	4+3-	20	50660694	4+3-	INS	-178	12	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50665426	2+2-	20	50665408	2+2-	INS	-111	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50666223	2+2-	20	50666228	2+2-	INS	-92	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50672395	4+5-	20	50672466	4+5-	ITX	-127	53	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50677238	3+1-	20	50677286	1+2-	INS	-201	35	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50680782	6+0-	20	50680910	0+3-	DEL	91	37	2	COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	50683918	2+3-	20	50683945	2+3-	INS	-108	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50691242	2+2-	20	50691383	2+3-	INS	-173	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50691496	2+1-	20	50691564	0+2-	INS	-211	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50699172	2+2-	20	50699148	2+2-	INS	-103	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50700029	2+0-	20	50700138	0+2-	INS	-206	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50701659	4+3-	20	50701749	4+3-	INS	-92	18	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50704773	2+2-	20	50704759	2+2-	INS	-108	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50710565	2+2-	20	50710573	2+2-	INS	-234	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50717714	3+3-	20	50717781	3+3-	INS	-274	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50726306	2+3-	20	50726333	2+3-	INS	-259	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50728407	2+2-	20	50728366	2+2-	INS	-97	38	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50745910	3+3-	20	50745924	3+3-	INS	-102	41	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50759449	2+0-	20	50759475	0+2-	INS	-310	28	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50770072	3+5-	20	50770239	3+5-	INS	-266	17	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50774742	2+0-	20	50774817	0+2-	INS	-254	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50785152	2+2-	20	50785172	2+2-	INS	-101	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50786357	2+3-	20	50786349	2+3-	INS	-117	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50791892	2+2-	20	50791866	2+2-	INS	-110	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50801051	2+4-	20	50801026	2+4-	INS	-116	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50809663	2+2-	20	50809660	2+2-	INS	-105	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50818029	3+0-	20	50818121	0+3-	INS	-188	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50852100	2+2-	20	50852066	2+2-	INS	-101	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50859299	2+0-	20	50859415	0+2-	INS	-208	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50862753	2+2-	20	50862718	2+2-	INS	-105	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50867720	2+0-	20	50867713	1+3-	INS	-255	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	50869359	2+2-	20	50869395	2+2-	INS	-108	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50880188	2+0-	20	50880267	0+2-	INS	-232	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50892325	2+2-	20	50892385	2+2-	INS	-98	25	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50904542	2+2-	20	50904590	2+2-	INS	-91	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50927827	2+2-	20	50927835	2+2-	INS	-224	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50944940	3+2-	20	50944954	3+2-	INS	-106	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50945477	2+2-	20	50945471	2+2-	INS	-243	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50946351	2+0-	20	50946379	2+2-	INS	-278	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50948861	2+0-	20	50949061	0+2-	INS	-115	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	50953444	3+5-	20	50953535	3+5-	INS	-153	25	3	COLO-829_v2_74|1:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	50965059	2+0-	20	50965067	0+2-	INS	-295	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	50981726	2+3-	20	50981786	2+3-	INS	-242	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51001766	3+2-	20	51001772	3+2-	INS	-385	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51007788	2+2-	20	51007770	2+2-	INS	-243	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51015617	2+0-	20	51015722	2+5-	INS	-148	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51028008	2+0-	20	51028120	0+3-	INS	-193	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51036659	2+3-	20	51036684	2+3-	INS	-96	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51037279	2+2-	20	51037234	2+2-	INS	-121	35	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51039485	3+5-	20	51039581	3+5-	INS	-285	23	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51041084	3+1-	20	51041400	36+72-	ITX	-160	99	36	COLO-829BL-IL|11:COLO-829-IL|25	0.30	BreakDancerMax-0.0.1r81	|q10|o20
20	51041382	32+1-	20	51041400	0+33-	DEL	154	99	31	COLO-829BL-IL|7:COLO-829-IL|24	0.26	BreakDancerMax-0.0.1r81	|q10|o20
20	51052748	2+3-	20	51052787	2+3-	INS	-100	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51068556	2+2-	20	51068541	2+2-	INS	-113	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51073311	2+1-	20	51073379	0+2-	INS	-241	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51084363	2+2-	20	51084380	1+2-	INS	-283	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51091008	3+1-	20	51091028	0+2-	INS	-241	35	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	51157137	2+1-	20	51157221	1+2-	INS	-218	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51170133	3+1-	20	51170274	0+2-	INS	-155	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51175361	2+2-	20	51175335	2+2-	INS	-106	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	51192547	2+0-	20	51192544	2+4-	INS	-263	34	4	COLO-829_v2_74|3:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	51202875	2+0-	20	51202879	0+2-	INS	-294	16	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	51216947	2+0-	20	51217024	2+2-	INS	-243	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51217133	2+0-	20	51217262	0+3-	INS	-203	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51224700	2+2-	20	51224662	2+2-	INS	-98	33	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	51246100	2+2-	20	51246076	2+2-	INS	-114	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51251188	2+2-	20	51251182	2+2-	INS	-91	27	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51254097	20+21-	20	51254079	20+21-	ITX	-144	99	12	COLO-829BL-IL|6:COLO-829-IL|6	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	51262081	2+2-	20	51262070	2+2-	INS	-108	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51275166	2+2-	20	51275176	2+2-	INS	-107	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51278586	2+0-	20	51278980	0+2-	DEL	80	52	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51288250	2+2-	20	51288242	2+2-	INS	-116	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51292666	2+3-	20	51292729	2+3-	INS	-108	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51303682	2+3-	20	51303665	2+3-	INS	-240	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51313228	2+2-	20	51313223	2+2-	INS	-102	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51314326	2+2-	20	51314311	2+2-	INS	-249	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51355652	3+3-	20	51355658	3+3-	INS	-112	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	51399278	3+3-	20	51399264	3+3-	INS	-108	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51401826	3+4-	20	51401839	3+4-	INS	-98	38	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51404814	3+3-	20	51404806	3+3-	INS	-279	33	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51414306	2+2-	20	51414272	2+2-	INS	-102	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	51416124	3+1-	20	51416192	1+2-	INS	-176	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	51426072	2+2-	20	51426040	2+2-	INS	-93	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51454038	2+2-	20	51454039	2+2-	INS	-217	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51457443	5+4-	20	51457500	5+4-	INS	-276	34	4	COLO-829_v2_74|3:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51465620	2+0-	20	51465607	24+27-	INS	-101	99	26	COLO-829BL-IL|8:COLO-829_v2_74|2:COLO-829-IL|16	0.37	BreakDancerMax-0.0.1r81	|q10|o20
20	51468834	2+3-	20	51468821	2+3-	INS	-250	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51473410	3+2-	20	51473369	3+2-	INS	-121	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51496913	3+3-	20	51496927	3+3-	INS	-253	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51519497	7+1-	20	51519713	2+5-	DEL	190	58	3	COLO-829-IL|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	51519497	4+1-	20	51519594	1+4-	DEL	112	53	3	COLO-829BL-IL|1:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	51532702	4+10-	20	51533149	2+11-	DEL	514	79	4	COLO-829BL-IL|4	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	51532702	0+10-	20	51532970	15+2-	ITX	131	99	9	COLO-829BL-IL|2:COLO-829-IL|7	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	51537513	2+2-	20	51537491	2+2-	INS	-96	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51537991	2+3-	20	51538004	2+3-	INS	-115	29	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51544355	2+1-	20	51544412	0+2-	INS	-250	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51553038	3+2-	20	51553037	3+2-	INS	-98	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51567090	3+2-	20	51567135	3+2-	INS	-233	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51568821	3+2-	20	51568857	3+2-	INS	-205	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51607034	2+0-	20	51607176	0+2-	INS	-185	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51607528	3+2-	20	51607510	3+2-	INS	-106	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51609074	4+3-	20	51609190	0+2-	INS	-180	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51618210	4+1-	20	51618239	0+3-	INS	-252	38	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	51682097	3+2-	20	51682082	3+2-	INS	-96	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51696350	3+1-	20	51696443	0+3-	INS	-192	38	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	51722732	2+0-	20	51722924	0+2-	INS	-138	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51728816	2+2-	20	51728765	2+2-	INS	-401	30	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51740804	2+3-	20	51740792	2+3-	INS	-99	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51757464	2+3-	20	51757485	2+3-	INS	-233	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51769107	4+0-	20	51769945	1+22-	DEL	582	72	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51769382	21+0-	20	51769945	1+19-	DEL	575	99	18	COLO-829BL-IL|9:COLO-829-IL|9	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	51780704	2+4-	20	51780728	2+4-	INS	-108	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51787102	2+2-	20	51787102	2+2-	INS	-104	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51794396	2+1-	20	51794530	0+3-	INS	-214	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51817377	2+4-	20	51817351	2+4-	INS	-409	23	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51820292	2+2-	20	51820269	2+2-	INS	-111	30	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51844590	6+6-	20	51849258	8+0-	INV	4572	99	6	COLO-829BL-IL|3:COLO-829-IL|3	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	51844590	0+6-	20	51849504	1+9-	INV	4866	99	6	COLO-829BL-IL|2:COLO-829-IL|4	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	51845119	2+2-	20	51845080	2+2-	INS	-104	37	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51845443	3+3-	20	51845496	3+3-	INS	-388	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51865803	2+2-	20	51865766	2+2-	INS	-99	37	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51884020	2+3-	20	51884000	2+3-	INS	-96	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51887615	52+44-	20	51887793	52+44-	INS	-98	99	35	COLO-829BL-IL|11:COLO-829-IL|24	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	51890488	2+0-	20	51890556	0+2-	INS	-239	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51891329	3+0-	20	51891826	0+3-	DEL	196	79	3	COLO-829_v2_74|3	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	51891438	6+0-	20	51891653	0+6-	DEL	181	99	6	COLO-829-IL|6	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	51897730	2+3-	20	51897728	2+3-	INS	-102	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51897934	3+3-	20	51897990	3+3-	INS	-112	33	3	COLO-829BL-IL|1:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	51911164	2+2-	20	51911164	2+2-	INS	-90	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51913118	2+2-	20	51913083	2+2-	INS	-110	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51913706	27+1-	20	51913735	0+28-	DEL	99	99	27	COLO-829BL-IL|14:COLO-829-IL|13	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	51915433	3+4-	20	51915481	3+4-	INS	-287	27	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51921916	3+0-	20	51922020	0+3-	INS	-222	33	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51956373	4+4-	20	51956529	4+4-	INS	-251	10	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51963211	4+4-	20	51963246	4+4-	INS	-90	50	4	COLO-829BL-IL|1:COLO-829-IL|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	51975303	2+3-	20	51975331	2+3-	INS	-98	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51981302	3+2-	20	51981282	3+2-	INS	-117	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51982655	3+2-	20	51982616	3+2-	INS	-114	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	51983240	2+2-	20	51983200	2+2-	INS	-116	34	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	51995617	2+3-	20	51995591	2+3-	INS	-111	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52022129	2+1-	20	52022234	1+3-	INS	-126	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52025702	2+2-	20	52025682	2+2-	INS	-387	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52032341	2+0-	20	52032478	1+3-	INS	-160	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52043480	2+0-	20	52043555	1+4-	INS	-168	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	52045302	3+3-	20	52045357	3+3-	INS	-168	32	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52046260	2+2-	20	52046250	2+2-	INS	-104	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52055247	3+3-	20	52055268	3+3-	INS	-93	37	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52070409	3+3-	20	52070413	3+3-	INS	-118	43	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52072262	2+0-	20	52072276	0+2-	INS	-265	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52076559	3+0-	20	52076590	0+2-	INS	-275	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52083639	3+0-	20	52083644	0+3-	INS	-214	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52094448	3+2-	20	52094488	3+2-	INS	-106	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52106223	2+2-	20	52106251	2+2-	INS	-100	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52107791	2+1-	20	52107865	1+3-	INS	-124	22	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52111797	2+2-	20	52111792	2+2-	INS	-84	31	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52131621	2+2-	20	52131623	2+2-	INS	-100	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52135042	2+2-	20	52135041	2+2-	INS	-229	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52140386	2+2-	20	52140378	2+2-	INS	-114	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52154536	2+2-	20	52154558	2+2-	INS	-108	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52156227	2+0-	20	52156208	0+2-	INS	-209	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52168842	2+0-	20	52168994	0+2-	INS	-160	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52191936	4+5-	20	52192043	4+5-	INS	-157	33	4	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52195305	2+2-	20	52195268	2+2-	INS	-116	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52200884	2+0-	20	52200909	0+2-	INS	-297	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52204474	2+0-	20	52204573	0+2-	INS	-221	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52215026	2+2-	20	52215053	2+2-	INS	-247	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52239629	2+2-	20	52239590	2+2-	INS	-98	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52252556	3+4-	20	52252591	3+4-	INS	-287	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52254889	2+4-	20	52254919	2+4-	INS	-93	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52277911	3+3-	20	52277918	3+3-	INS	-195	32	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52295768	2+2-	20	52295766	2+2-	INS	-106	27	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52332018	2+2-	20	52331997	2+2-	INS	-112	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52342405	3+3-	20	52342489	3+3-	INS	-105	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52350236	2+3-	20	52350263	2+3-	INS	-89	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52353665	2+2-	20	52353716	2+2-	INS	-340	15	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52371995	2+3-	20	52372024	2+3-	INS	-106	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52374332	3+1-	20	52374474	2+4-	INS	-116	36	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52375412	2+2-	20	52375394	2+2-	INS	-107	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52376123	2+3-	20	52376111	2+3-	INS	-98	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52379356	2+2-	20	52379325	2+2-	INS	-101	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52388478	3+2-	20	52388440	3+2-	INS	-250	28	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52389129	3+3-	20	52389193	3+3-	INS	-192	25	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52396277	2+0-	20	52396465	1+2-	INS	-115	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52402112	3+3-	20	52402249	2+2-	INS	-151	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52404495	2+3-	20	52404480	2+3-	INS	-107	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52408937	3+3-	20	52408960	3+3-	INS	-251	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52417974	2+0-	20	52418129	0+2-	INS	-156	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52418076	2+2-	20	52418045	2+2-	INS	-105	36	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52437205	3+2-	20	52437206	0+3-	INS	-238	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	52470646	3+1-	20	52470789	1+2-	INS	-144	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52475586	2+2-	20	52475582	2+2-	INS	-106	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52476059	5+4-	20	52476081	5+4-	INS	-104	37	3	COLO-829BL-IL|1:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	52504681	4+1-	20	52504691	0+3-	INS	-242	39	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	52509158	2+2-	20	52509143	2+2-	INS	-104	33	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52521399	3+1-	20	52521454	1+3-	INS	-212	27	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	52533186	2+2-	20	52533153	2+2-	INS	-106	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52548774	2+2-	20	52548782	2+2-	INS	-247	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52551593	2+3-	20	52551583	2+3-	INS	-105	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52558310	3+3-	20	52558347	3+3-	INS	-105	27	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52559712	2+2-	20	52559723	2+2-	INS	-103	29	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52584138	2+2-	20	52584122	2+2-	INS	-106	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52591121	3+0-	20	52591188	0+3-	INS	-274	46	3	COLO-829_v2_74|3	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	52607330	2+2-	20	52607319	2+2-	INS	-111	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52616467	2+1-	20	52616548	0+4-	INS	-183	18	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	52628902	2+2-	20	52628898	2+2-	INS	-100	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52636062	2+4-	20	52636132	2+4-	INS	-93	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52638684	3+3-	20	52638703	3+3-	ITX	-128	38	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52650607	3+2-	20	52650640	3+2-	INS	-348	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52668739	2+2-	20	52668703	2+2-	INS	-385	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52683400	2+2-	20	52683505	2+4-	INS	-295	40	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52695292	2+0-	20	52695423	0+2-	DEL	85	49	2	COLO-829-IL|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	52700152	2+0-	20	52700203	0+3-	INS	-259	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52702314	2+1-	20	52702387	0+2-	INS	-240	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52723214	2+2-	20	52723167	2+2-	INS	-114	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52725781	5+0-	20	52726368	1+94-	DEL	320	99	5	COLO-829_v2_74|5	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	52726131	89+2-	20	52726368	0+88-	DEL	318	99	88	COLO-829BL-IL|23:COLO-829_v2_74|16:COLO-829-IL|49	0.44	BreakDancerMax-0.0.1r81	|q10|o20
20	52737515	3+4-	20	52737485	3+4-	INS	-108	50	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52738718	4+2-	20	52738779	1+2-	INS	-188	24	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52742037	2+3-	20	52742072	2+3-	INS	-226	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52745819	2+2-	20	52745797	2+2-	INS	-96	34	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52756364	2+2-	20	52756311	2+2-	INS	-403	31	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52762092	2+2-	20	52762121	2+2-	INS	-243	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52774700	2+2-	20	52774692	2+2-	INS	-112	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52792431	2+2-	20	52792404	2+2-	INS	-111	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52794998	3+3-	20	52795048	3+3-	INS	-103	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52811481	3+3-	20	52811610	3+3-	INS	-213	19	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52825545	2+2-	20	52825497	2+2-	INS	-397	29	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52839335	2+2-	20	52839333	2+2-	INS	-90	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52849417	2+2-	20	52849449	2+2-	INS	-227	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52869053	1+5-	20	52869669	0+4-	INV	530	99	4	COLO-829BL-IL|1:COLO-829-IL|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	52881082	2+2-	20	52881096	2+2-	INS	-101	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	52888337	4+2-	20	52888408	4+2-	INS	-106	25	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52900084	2+4-	20	52900111	0+2-	INS	-310	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52913223	2+2-	20	52913187	2+2-	INS	-385	25	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52927309	2+2-	20	52927346	2+2-	INS	-214	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	52944329	2+2-	20	52944331	2+2-	INS	-89	26	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	52978212	2+2-	20	52978166	2+2-	INS	-119	36	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	52982170	3+3-	20	52982213	3+3-	INS	-109	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53012988	2+0-	20	53013023	1+3-	INS	-235	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	53014535	3+2-	20	53014614	3+2-	INS	-100	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53022300	3+3-	20	53022294	3+3-	INS	-108	27	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53037915	2+2-	20	53037897	2+2-	INS	-112	33	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53051298	2+2-	20	53051267	2+2-	INS	-398	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53054924	2+4-	20	53054974	2+4-	INS	-102	26	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53056664	2+2-	20	53056643	2+2-	INS	-112	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53071300	2+2-	20	53071266	2+2-	INS	-98	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53077354	2+2-	20	53077363	2+2-	INS	-102	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53104647	2+2-	20	53104619	2+2-	INS	-104	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53122329	2+2-	20	53122320	2+2-	INS	-106	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53143097	2+2-	20	53143109	2+2-	INS	-106	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53145243	2+1-	20	53145319	1+2-	INS	-273	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53146665	2+0-	20	53146803	0+2-	INS	-176	15	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	53169143	3+3-	20	53169183	3+3-	INS	-164	28	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53175205	2+2-	20	53175164	2+2-	INS	-122	34	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53179538	2+1-	20	53179640	2+2-	INS	-136	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53179791	2+0-	20	53179930	0+2-	INS	-142	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53182819	2+2-	20	53182848	2+2-	INS	-211	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53195319	2+9-	20	53195342	2+9-	INS	-90	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53197384	2+2-	20	53197353	2+2-	INS	-97	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53198236	2+0-	20	53198343	1+3-	INS	-157	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53199046	2+1-	20	53199235	2+2-	INS	-118	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53199371	2+0-	20	53199466	1+2-	INS	-202	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53205643	3+0-	20	53205760	0+3-	INS	-203	34	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	53225507	2+2-	20	53225452	2+2-	INS	-404	32	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53240611	3+2-	20	53240620	3+2-	INS	-88	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53261648	3+3-	20	53261690	3+3-	INS	-192	28	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53311619	2+0-	20	53311697	0+2-	INS	-249	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53330224	2+1-	20	53330242	0+2-	INS	-330	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53332688	3+3-	20	53332702	3+3-	INS	-186	31	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53342395	2+2-	20	53342384	2+2-	INS	-104	32	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53351626	2+0-	20	53351701	0+2-	INS	-245	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53372290	3+2-	20	53372277	3+2-	INS	-100	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53380783	2+2-	20	53380784	2+2-	INS	-105	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53388349	3+1-	20	53388436	0+2-	INS	-184	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53393015	3+4-	20	53393029	3+4-	INS	-299	29	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53397262	46+0-	20	53397554	3+7-	DEL	92	90	4	COLO-829_v2_74|4	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	53397262	42+0-	20	53397287	0+45-	DEL	96	99	42	COLO-829BL-IL|12:COLO-829-IL|30	0.38	BreakDancerMax-0.0.1r81	|q10|o20
20	53399788	2+2-	20	53399740	2+2-	INS	-111	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53413571	2+0-	20	53413691	0+2-	INS	-210	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53427915	2+3-	20	53427993	2+3-	INS	-99	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53473850	2+0-	20	53473955	0+3-	INS	-200	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53476751	2+2-	20	53476714	2+2-	INS	-95	37	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53486317	2+2-	20	53486260	2+2-	ITX	-130	54	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53493080	2+3-	20	53493091	2+3-	INS	-95	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53507105	5+2-	20	53507165	5+2-	INS	-99	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53507235	3+0-	20	53507379	0+3-	INS	-167	22	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53517292	3+3-	20	53517315	3+3-	INS	-107	37	3	COLO-829BL-IL|1:COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53535883	2+0-	20	53535976	1+3-	INS	-168	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53544267	2+2-	20	53544260	2+2-	INS	-95	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53546663	2+2-	20	53546648	2+2-	INS	-107	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53547637	29+8-	20	53547912	5+21-	DEL	329	99	17	COLO-829BL-IL|5:COLO-829-IL|12	1.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53558896	2+3-	20	53558959	2+3-	INS	-101	25	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53571233	3+2-	20	53571223	3+2-	INS	-95	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53576395	2+3-	20	53576376	2+3-	INS	-231	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53590870	2+2-	20	53590868	2+2-	INS	-101	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53613865	2+2-	20	53613838	2+2-	INS	-99	35	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53618363	2+2-	20	53618324	2+2-	INS	-105	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53621282	6+5-	20	53621497	6+5-	INS	-94	19	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53640957	2+2-	20	53640977	2+2-	INS	-88	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53644597	3+2-	20	53644632	3+2-	INS	-388	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53644832	3+0-	20	53645009	1+4-	INS	-104	38	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	53650617	3+3-	20	53650615	3+3-	INS	-115	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53657979	2+2-	20	53657953	2+2-	INS	-250	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53674645	3+2-	20	53674626	3+2-	INS	-104	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53684572	2+2-	20	53684578	2+2-	INS	-107	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53696919	3+4-	20	53696899	3+4-	INS	-95	29	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53719369	2+3-	20	53719383	2+3-	INS	-102	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53741586	2+3-	20	53741598	2+3-	INS	-226	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53749077	3+2-	20	53749139	3+2-	INS	-324	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53749514	3+2-	20	53749604	3+2-	INS	-175	13	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53773359	4+3-	20	53773390	4+3-	INS	-211	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53774373	2+2-	20	53774353	2+2-	INS	-88	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53779695	3+3-	20	53779753	3+3-	INS	-378	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53796610	2+2-	20	53796622	2+2-	INS	-87	29	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53802178	3+3-	20	53802201	3+3-	ITX	-127	37	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53807837	2+3-	20	53807886	2+3-	INS	-103	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53819286	2+0-	20	53819442	0+2-	INS	-165	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53825054	3+2-	20	53825036	3+2-	INS	-110	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53835850	2+2-	20	53835821	2+2-	INS	-236	26	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53840085	24+23-	20	53840090	24+23-	INS	-101	99	19	COLO-829BL-IL|5:COLO-829-IL|14	0.23	BreakDancerMax-0.0.1r81	|q10|o20
20	53851837	2+2-	20	53851805	2+2-	INS	-103	32	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53853062	3+3-	20	53853135	3+3-	INS	-88	25	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53860182	2+0-	20	53860287	0+2-	INS	-210	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53867789	2+2-	20	53874017	1+36-	DEL	5996	44	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53868054	38+0-	20	53874017	1+34-	DEL	6004	99	32	COLO-829BL-IL|8:COLO-829_v2_74|1:COLO-829-IL|23	0.48	BreakDancerMax-0.0.1r81	|q10|o20
20	53868054	6+0-	20	53874253	1+9-	DEL	5992	99	6	COLO-829_v2_74|6	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	53884339	2+3-	20	53884313	2+3-	INS	-251	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53885023	2+2-	20	53885011	2+2-	INS	-239	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	53896003	2+1-	20	53896008	3+3-	INS	-149	25	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	53896178	2+0-	20	53896262	0+2-	INS	-191	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53896642	59+0-	20	53896941	0+49-	DEL	319	99	48	COLO-829BL-IL|17:COLO-829-IL|31	0.42	BreakDancerMax-0.0.1r81	|q10|o20
20	53896642	11+0-	20	53897068	4+13-	DEL	324	99	11	COLO-829_v2_74|11	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	53897467	3+1-	20	53897548	0+2-	INS	-249	7	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53902372	2+1-	20	53902456	1+2-	INS	-246	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53903079	2+2-	20	53903068	2+2-	INS	-111	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53912937	6+5-	20	53912993	6+5-	INS	-98	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	53920309	4+1-	20	53920394	0+4-	DEL	92	75	4	COLO-829BL-IL|1:COLO-829-IL|3	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	53924573	3+6-	20	53924635	3+6-	INS	-112	35	3	COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53953955	12+0-	20	53953995	0+12-	DEL	90	99	12	COLO-829BL-IL|2:COLO-829-IL|10	0.28	BreakDancerMax-0.0.1r81	|q10|o20
20	53955126	2+0-	20	53955130	1+3-	INS	-229	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	53961396	2+2-	20	53961369	2+2-	INS	-106	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53975816	8+6-	20	53976054	2+7-	INS	-98	75	6	COLO-829BL-IL|3:COLO-829-IL|3	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	53976214	2+5-	20	53976199	0+3-	INS	-364	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	53975950	5+0-	20	53976054	0+5-	DEL	89	96	5	COLO-829BL-IL|2:COLO-829-IL|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	53978020	2+2-	20	53978046	2+2-	INS	-212	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	53997955	2+2-	20	53997925	2+2-	INS	-112	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54002708	2+2-	20	54002702	2+2-	INS	-104	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54010201	2+3-	20	54010224	2+3-	INS	-230	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54021422	4+3-	20	54021504	4+3-	INS	-101	34	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54043492	2+0-	20	54043561	1+3-	INS	-164	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54050138	2+3-	20	54050214	2+3-	INS	-91	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54056351	2+0-	20	54056348	0+2-	INS	-218	27	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	54078065	3+2-	20	54078083	3+2-	INS	-110	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54081147	2+0-	20	54081304	1+2-	INS	-160	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54084052	2+2-	20	54084086	2+2-	INS	-93	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	54086619	4+0-	20	54086684	0+4-	INS	-221	31	4	COLO-829_v2_74|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	54088446	2+2-	20	54088502	2+2-	INS	-247	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54096504	2+3-	20	54096527	2+3-	INS	-376	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54111001	2+2-	20	54111041	2+2-	INS	-236	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	54127174	2+2-	20	54127152	2+2-	INS	-371	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54135050	3+3-	20	54135100	3+3-	INS	-169	27	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54138502	2+0-	20	54138576	1+3-	INS	-196	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54144535	3+3-	20	54144532	3+3-	INS	-107	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54153317	2+2-	20	54153281	2+2-	INS	-98	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54162673	2+0-	20	54162831	0+2-	INS	-149	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54209147	2+1-	20	54209305	0+2-	INS	-181	26	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	54216525	2+2-	20	54216598	1+3-	INS	-132	23	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54264420	3+1-	20	54264531	2+2-	INS	-128	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54264995	3+2-	20	54265058	3+2-	INS	-215	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54292817	7+0-	20	54292798	0+7-	INS	-94	99	7	COLO-829BL-IL|2:COLO-829-IL|5	0.17	BreakDancerMax-0.0.1r81	|q10|o20
20	54297880	2+3-	20	54297915	2+3-	INS	-113	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54310332	3+3-	20	54310378	3+3-	INS	-198	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54320791	3+3-	20	54320743	3+3-	INS	-112	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54344652	3+3-	20	54344725	3+3-	INS	-90	25	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54381710	3+2-	20	54381772	3+2-	INS	-187	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	54391500	2+2-	20	54391507	2+2-	INS	-99	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54394566	3+3-	20	54394648	3+3-	INS	-91	19	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54434989	2+2-	20	54435023	2+2-	INS	-245	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54462690	4+4-	20	54462691	4+4-	INS	-236	50	4	COLO-829BL-IL|2:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54472682	2+3-	20	54472670	2+3-	INS	-95	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54475990	3+1-	20	54476023	0+2-	INS	-199	28	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	54505440	2+0-	20	54505466	1+3-	INS	-302	25	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54518085	3+3-	20	54518127	3+3-	INS	-102	27	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54525717	2+3-	20	54525728	2+3-	INS	-339	18	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	54534894	11+0-	20	54545271	5+11-	DEL	10377	99	11	COLO-829BL-IL|4:COLO-829-IL|7	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	54535113	0+5-	20	54545271	5+0-	ITX	9974	99	5	COLO-829BL-IL|4:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54535642	2+0-	20	54535843	0+2-	INS	-120	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54537226	3+3-	20	54537265	1+2-	INS	-218	27	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54566947	2+2-	20	54566968	2+2-	INS	-107	24	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54574260	2+3-	20	54574272	2+3-	INS	-97	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54585159	2+2-	20	54585167	2+2-	INS	-101	30	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	54632732	3+3-	20	54632788	3+3-	INS	-102	35	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54661954	2+2-	20	54661980	2+2-	INS	-99	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	54694898	2+2-	20	54694865	2+2-	INS	-116	36	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54699407	2+2-	20	54699369	2+2-	INS	-387	26	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54719300	12+11-	20	54719386	12+11-	ITX	-196	99	8	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|5	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	54732854	2+2-	20	54732835	2+2-	INS	-93	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54734714	4+2-	20	54734752	4+2-	INS	-125	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54746198	2+1-	20	54746196	0+2-	INS	-293	19	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	54758482	2+0-	20	54758487	2+3-	INS	-223	24	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	54770983	2+2-	20	54771016	2+2-	INS	-247	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54771560	2+2-	20	54771511	2+2-	INS	-259	32	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	54774778	0+2-	20	54775949	0+3-	INV	1059	58	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54778529	3+0-	20	54778684	0+3-	INS	-163	37	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54786062	2+2-	20	54786031	2+2-	INS	-381	24	2	COLO-829_v2_74|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	54796256	3+3-	20	54796323	3+3-	INS	-241	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	54807453	4+1-	20	54807486	1+2-	INS	-295	32	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54808391	3+1-	20	54808503	1+3-	INS	-156	42	4	COLO-829_v2_74|2:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54814196	2+0-	20	54814296	0+2-	INS	-222	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54816332	2+0-	20	54816511	0+2-	INS	-147	23	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	54836512	2+3-	20	54836479	2+3-	INS	-125	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54839590	3+3-	20	54839610	3+3-	INS	-402	17	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	54840469	2+3-	20	54840441	2+3-	INS	-105	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54864540	2+2-	20	54864496	2+2-	INS	-109	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	54901708	2+2-	20	54901690	2+2-	INS	-115	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	54906339	2+0-	20	54906372	1+3-	INS	-225	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	54909495	2+2-	20	54909462	2+2-	INS	-383	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54930584	3+0-	20	54930701	0+2-	INS	-187	17	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	54935944	2+2-	20	54935938	2+2-	INS	-111	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54945425	2+2-	20	54945450	2+2-	INS	-103	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54954794	3+3-	20	54954802	3+3-	INS	-266	30	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	54957048	2+2-	20	54957050	3+3-	INS	-189	20	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	54957777	2+3-	20	54957758	2+3-	INS	-98	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54972496	3+4-	20	54972587	3+4-	INS	-105	24	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	54981359	2+4-	20	54981400	2+4-	INS	-357	16	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55003229	2+2-	20	55003187	2+2-	INS	-392	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55022214	2+2-	20	55022169	2+2-	INS	-104	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55023654	3+0-	20	55023669	1+4-	INS	-238	13	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55032754	2+2-	20	55032759	2+2-	INS	-113	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55040407	57+2-	20	55040423	1+44-	DEL	108	99	43	COLO-829BL-IL|17:COLO-829-IL|26	0.16	BreakDancerMax-0.0.1r81	|q10|o20
20	55040407	14+2-	20	55040611	0+9-	DEL	107	99	8	COLO-829_v2_74|8	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	55064319	2+2-	20	55064328	2+2-	INS	-103	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55070195	2+1-	20	55070366	1+3-	INS	-155	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55075122	2+0-	20	55075116	0+2-	INS	-285	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55090072	3+2-	20	55090144	0+2-	INS	-194	18	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55099580	8+2-	20	55099684	0+5-	INS	-149	33	4	COLO-829_v2_74|4	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	55099580	2+1-	20	55099578	2+2-	DEL	92	33	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	55106208	3+2-	20	55106246	3+2-	INS	-93	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55118966	14+1-	20	55119058	0+10-	DEL	126	99	10	COLO-829BL-IL|4:COLO-829-IL|6	0.33	BreakDancerMax-0.0.1r81	|q10|o20
20	55118966	3+0-	20	55119369	0+3-	DEL	140	46	2	COLO-829_v2_74|2	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	55120082	2+1-	20	55120170	0+2-	INS	-243	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55133257	2+2-	20	55133242	2+2-	INS	-92	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55135023	4+6-	20	55135102	4+6-	INS	-110	48	4	COLO-829-IL|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55135952	2+2-	20	55135956	2+2-	INS	-100	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55162267	2+3-	20	55162277	2+3-	INS	-101	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55184414	4+3-	20	55184444	0+2-	INS	-174	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55198621	4+0-	20	55198901	0+16-	DEL	89	92	4	COLO-829_v2_74|4	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	55198882	14+0-	20	55198901	0+12-	DEL	94	99	11	COLO-829BL-IL|2:COLO-829-IL|9	0.23	BreakDancerMax-0.0.1r81	|q10|o20
20	55198882	3+0-	20	55199266	0+3-	DEL	79	71	3	COLO-829_v2_74|3	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	55212883	2+2-	20	55212900	2+2-	INS	-100	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55227052	7+7-	20	55227439	4+4-	ITX	201	43	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55240959	3+4-	20	55241022	3+4-	INS	-159	25	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55245648	2+3-	20	55245655	2+3-	INS	-214	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55254770	2+0-	20	55254886	1+2-	INS	-183	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55293214	2+3-	20	55293248	2+3-	INS	-95	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55305182	2+2-	20	55305160	2+2-	INS	-231	25	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55312689	3+0-	20	55312883	0+3-	INS	-140	35	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	55341474	4+0-	20	55341543	3+2-	INS	-278	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55341678	3+0-	20	55341694	0+4-	INS	-230	22	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	55346073	2+2-	20	55346093	2+2-	INS	-103	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55358361	2+3-	20	55358373	2+3-	INS	-102	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55377228	2+2-	20	55377224	2+2-	INS	-239	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55387100	2+2-	20	55387134	2+2-	INS	-94	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55387374	2+3-	20	55387421	2+3-	INS	-235	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55425769	10+1-	20	55425805	27+26-	INS	-119	99	23	COLO-829BL-IL|4:COLO-829_v2_74|9:COLO-829-IL|10	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	55426064	10+0-	20	55426050	0+10-	INS	-126	77	10	COLO-829_v2_74|8:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	55426543	2+2-	20	55426526	2+2-	INS	-104	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55470597	3+5-	20	55470667	3+5-	INS	-327	24	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55473469	3+3-	20	55473519	3+3-	INS	-103	22	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55473658	2+2-	20	55473635	2+2-	INS	-373	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55483768	2+2-	20	55483733	2+2-	INS	-90	36	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55498509	3+3-	20	55498548	3+3-	INS	-107	23	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	55515281	2+2-	20	55515281	2+2-	INS	-100	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55521243	3+3-	20	55521254	3+3-	INS	-291	31	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55529628	2+0-	20	55529830	0+2-	INS	-124	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55531046	3+0-	20	55531051	0+2-	INS	-169	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55568780	2+2-	20	55568780	2+2-	INS	-220	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55576042	2+0-	20	55576088	0+2-	INS	-278	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55580335	2+3-	20	55580320	2+3-	INS	-104	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55583677	2+3-	20	55583646	2+3-	INS	-110	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55585945	2+2-	20	55585950	2+2-	INS	-98	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55587738	6+2-	20	55587784	8+14-	INS	-99	99	9	COLO-829BL-IL|3:COLO-829-IL|6	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	55594263	2+2-	20	55594306	2+2-	INS	-195	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55596290	2+0-	20	55596405	0+2-	INS	-217	25	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55596738	2+2-	20	55596731	2+2-	INS	-93	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55621006	2+2-	20	55620994	2+2-	INS	-100	32	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55621742	4+4-	20	55621748	4+4-	INS	-251	45	4	COLO-829_v2_74|2:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55640276	2+2-	20	55640249	2+2-	INS	-376	23	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55646832	3+4-	20	55646906	3+4-	INS	-233	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55668983	2+0-	20	55669093	1+2-	INS	-226	27	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55696841	3+1-	20	55697018	0+2-	INS	-122	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55704219	2+0-	20	55704357	0+2-	INS	-193	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55742059	2+0-	20	55742112	1+3-	INS	-175	27	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	55766223	2+2-	20	55766165	2+2-	INS	-408	34	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	55767548	5+3-	20	55767681	5+3-	INS	-136	26	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55769383	2+3-	20	55769351	2+3-	INS	-255	25	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	55789754	2+2-	20	55789745	1+4-	INS	-202	23	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55794324	2+2-	20	55794312	2+2-	INS	-240	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55807202	2+2-	20	55807227	2+2-	INS	-237	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55824550	3+2-	20	55824564	3+2-	INS	-230	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55847898	2+2-	20	55847900	2+2-	INS	-104	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55854894	2+2-	20	55854909	2+2-	INS	-94	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55865162	2+2-	20	55865190	2+2-	INS	-107	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55870022	2+1-	20	55870172	0+2-	INS	-157	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55896900	3+1-	20	55896893	0+3-	INS	-195	20	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55923015	3+1-	20	55923009	0+2-	INS	-238	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55939735	2+3-	20	55939776	2+3-	INS	-203	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55951229	6+4-	20	55951347	6+4-	INS	-285	19	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55951417	3+1-	20	55951442	0+2-	INS	-300	11	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55957432	7+3-	20	55957427	9+0-	ITX	-149	53	3	COLO-829BL-IL|1:COLO-829-IL|2	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	55957432	7+0-	20	55957788	0+16-	DEL	305	99	6	COLO-829BL-IL|4:COLO-829_v2_74|1:COLO-829-IL|1	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	55957572	6+0-	20	55957906	0+2-	DEL	362	36	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	55957572	4+0-	20	55957788	0+10-	DEL	170	35	2	COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	55957572	2+0-	20	55957693	0+2-	DEL	91	42	2	COLO-829BL-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	55957706	8+0-	20	55957788	0+8-	DEL	92	99	8	COLO-829BL-IL|2:COLO-829-IL|6	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	55966275	2+0-	20	55966307	3+5-	INS	-178	43	4	COLO-829BL-IL|2:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	55971115	2+2-	20	55971106	2+2-	INS	-359	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55975229	2+2-	20	55975233	2+2-	INS	-103	30	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	55979042	2+0-	20	55979119	0+2-	INS	-257	26	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	55983358	11+0-	20	55983360	1+10-	DEL	89	99	7	COLO-829BL-IL|1:COLO-829-IL|6	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	55985663	4+2-	20	55985751	0+3-	INS	-181	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	55987996	26+0-	20	55988062	0+24-	DEL	106	99	22	COLO-829BL-IL|8:COLO-829-IL|14	0.20	BreakDancerMax-0.0.1r81	|q10|o20
20	55987996	3+0-	20	55988316	0+3-	DEL	102	68	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	56006165	2+1-	20	56006184	0+2-	INS	-308	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56026893	2+2-	20	56026892	2+2-	INS	-110	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56037091	2+0-	20	56037296	0+2-	INS	-120	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56037472	2+2-	20	56037503	2+2-	INS	-329	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56037982	3+2-	20	56037991	3+2-	INS	-101	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56040341	2+0-	20	56040391	0+2-	INS	-273	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56049972	3+3-	20	56049992	3+3-	INS	-103	40	3	COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56061507	2+4-	20	56061558	2+4-	INS	-113	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56064630	2+2-	20	56064773	0+2-	INS	-180	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56088882	2+2-	20	56088836	2+2-	INS	-111	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	56091082	2+2-	20	56091072	2+2-	INS	-106	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56094541	2+2-	20	56094566	2+2-	INS	-91	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	56105964	52+48-	20	56106040	0+4-	DEL	106	99	19	COLO-829BL-IL|8:COLO-829_v2_74|4:COLO-829-IL|7	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	56107789	2+3-	20	56107762	2+3-	INS	-111	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56120095	2+4-	20	56120133	2+4-	INS	-121	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56138770	2+0-	20	56138851	0+2-	INS	-233	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56149255	2+1-	20	56149264	0+2-	INS	-322	23	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	56151154	2+3-	20	56151134	2+3-	INS	-113	29	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	56157185	2+2-	20	56157160	2+2-	INS	-112	30	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	56171092	2+2-	20	56171058	2+2-	INS	-384	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56178499	2+2-	20	56178498	2+2-	INS	-94	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56201769	2+0-	20	56201867	0+2-	INS	-244	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56205106	38+43-	20	56205483	38+43-	INS	-99	99	13	COLO-829BL-IL|5:COLO-829-IL|8	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56208063	2+2-	20	56208054	2+2-	INS	-372	21	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	56237690	2+2-	20	56237663	2+2-	INS	-116	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56278955	2+2-	20	56278907	2+2-	INS	-111	40	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56282017	3+2-	20	56282012	3+2-	INS	-98	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56288985	3+3-	20	56289022	3+3-	INS	-272	26	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56294005	2+0-	20	56294128	1+2-	INS	-187	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56298838	2+2-	20	56298827	2+2-	INS	-115	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56300073	3+0-	20	56300067	6+3-	INS	-305	25	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	56308965	2+2-	20	56308976	2+2-	INS	-106	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56313692	3+1-	20	56313691	1+3-	INS	-189	34	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	56319541	3+4-	20	56319598	3+4-	INS	-160	26	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56337438	2+2-	20	56337419	2+2-	INS	-117	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56376968	2+3-	20	56377022	2+3-	INS	-251	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56403305	2+3-	20	56403317	2+3-	INS	-102	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56408112	3+2-	20	56408175	3+2-	INS	-330	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56417916	2+2-	20	56417874	2+2-	INS	-257	27	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56428209	2+2-	20	56428169	2+2-	INS	-109	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56433943	2+2-	20	56433913	2+2-	INS	-95	35	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56441147	2+2-	20	56441134	2+2-	INS	-108	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	56456705	2+2-	20	56456681	2+2-	INS	-103	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56479857	3+2-	20	56479898	3+2-	INS	-259	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56485647	2+3-	20	56485688	2+3-	INS	-225	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56491044	2+2-	20	56491029	2+2-	ITX	-132	43	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	56507330	3+3-	20	56507345	3+3-	INS	-187	31	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56524409	2+0-	20	56524586	1+2-	INS	-159	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56528628	19+19-	20	56528805	19+19-	INS	-94	99	17	COLO-829BL-IL|6:COLO-829-IL|11	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	56548020	2+3-	20	56548014	2+3-	INS	-90	31	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56550764	20+0-	20	56550867	0+22-	DEL	155	99	19	COLO-829BL-IL|11:COLO-829-IL|8	0.73	BreakDancerMax-0.0.1r81	|q10|o20
20	56568870	2+2-	20	56568890	2+2-	INS	-102	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	56573693	5+3-	20	56573800	5+3-	INS	-182	12	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56574027	2+2-	20	56573997	2+2-	INS	-91	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56585588	2+2-	20	56585586	2+2-	INS	-96	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56598161	2+0-	20	56598270	0+2-	INS	-173	18	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	56614728	2+2-	20	56614699	2+2-	INS	-378	24	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56622462	3+1-	20	56622645	0+2-	INS	-225	33	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56623925	2+2-	20	56624061	1+3-	INS	-144	20	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56628158	2+0-	20	56628242	1+3-	INS	-181	33	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56660412	2+2-	20	56660368	2+2-	INS	-258	28	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56661917	3+0-	20	56661902	0+2-	INS	-324	21	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	56663858	4+2-	20	56663932	4+2-	INS	-204	14	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56664002	2+0-	20	56664203	2+3-	INS	-138	18	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56676416	3+3-	20	56676436	3+3-	INS	-232	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56689355	3+1-	20	56689455	1+3-	INS	-239	26	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56699732	2+2-	20	56699734	2+2-	INS	-227	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56703319	5+0-	20	56703693	21+18-	INS	-380	66	7	COLO-829_v2_74|7	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	56703711	8+15-	20	56703693	12+5-	ITX	-332	99	9	COLO-829_v2_74|9	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56703862	3+1-	20	56703891	0+3-	INS	-224	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56705665	3+4-	20	56705674	3+4-	INS	-237	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56718138	2+0-	20	56718307	2+4-	INS	-131	39	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56732538	2+2-	20	56732582	2+2-	INS	-119	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56732783	2+2-	20	56732791	2+2-	INS	-102	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56755204	2+0-	20	56755270	0+2-	INS	-258	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56762949	2+2-	20	56762947	2+2-	INS	-241	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56572473	10+0-	20	56778559	1+74-	DEL	206118	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56783035	2+2-	20	56782998	2+2-	INS	-114	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56786193	2+0-	20	56786384	0+2-	INS	-134	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56791768	2+3-	20	56791729	2+3-	INS	-106	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56797314	2+2-	20	56797347	0+2-	INS	-174	11	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56814859	2+3-	20	56814843	2+3-	INS	-104	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	56816371	2+2-	20	56816327	2+2-	INS	-394	28	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	56822462	3+0-	20	56822481	0+3-	INS	-306	37	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	56822876	2+2-	20	56822878	2+2-	INS	-97	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56838951	12+1-	20	56839292	1+5-	DEL	130	67	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	56838951	8+0-	20	56839015	1+6-	DEL	91	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56878805	2+3-	20	56878831	2+3-	INS	-350	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56885912	2+2-	20	56885925	2+2-	ITX	-129	39	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56895305	2+2-	20	56895297	2+2-	INS	-394	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56913845	2+2-	20	56913836	2+2-	INS	-245	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56930783	3+3-	20	56930813	3+3-	INS	-243	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56936364	2+0-	20	56936514	0+2-	INS	-156	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56940408	3+2-	20	56940400	3+2-	INS	-392	20	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	56947895	3+3-	20	56947935	3+3-	INS	-104	37	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	56958756	2+0-	20	56958865	0+2-	INS	-212	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56963890	2+2-	20	56963888	2+2-	INS	-109	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56992222	2+3-	20	56992266	2+3-	INS	-221	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	56999364	2+2-	20	56999310	2+2-	INS	-404	32	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57044520	2+3-	20	57044541	2+3-	INS	-100	28	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57056792	3+2-	20	57056941	0+2-	INS	-137	33	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57071161	2+2-	20	57071198	2+2-	INS	-207	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57095352	2+2-	20	57095390	2+2-	INS	-87	27	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57114950	2+0-	20	57114938	1+3-	INS	-214	29	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	57131581	2+2-	20	57131585	2+2-	INS	-226	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57133777	2+2-	20	57133728	2+2-	INS	-399	29	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57137716	4+2-	20	57137744	4+2-	INS	-105	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57141607	12+3-	20	57141723	12+19-	DEL	95	99	11	COLO-829BL-IL|5:COLO-829-IL|6	0.30	BreakDancerMax-0.0.1r81	|q10|o20
20	57172974	3+0-	20	57173006	0+3-	INS	-221	23	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	57175288	3+0-	20	57175381	0+3-	INS	-217	34	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57182364	2+2-	20	57182350	2+2-	INS	-123	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57195066	2+0-	20	57195174	0+2-	INS	-209	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57197182	5+5-	20	57197295	5+5-	INS	-187	22	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57206320	4+4-	20	57206412	4+4-	INS	-158	23	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57208523	2+2-	20	57208563	2+2-	INS	-210	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57211623	2+2-	20	57211594	2+2-	INS	-107	31	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57219375	33+4-	20	57219505	1+31-	DEL	219	99	29	COLO-829BL-IL|11:COLO-829-IL|18	0.22	BreakDancerMax-0.0.1r81	|q10|o20
20	57219375	4+4-	20	57219684	0+6-	DEL	209	83	4	COLO-829_v2_74|4	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	57234263	2+2-	20	57234271	2+2-	INS	-219	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57250381	3+3-	20	57250381	3+3-	INS	-358	32	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57260236	2+3-	20	57260243	2+3-	INS	-112	26	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57269659	2+2-	20	57269651	2+2-	INS	-243	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57277483	4+1-	20	57277488	0+3-	INS	-199	35	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	57292633	2+2-	20	57292615	2+2-	INS	-368	22	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57293413	2+2-	20	57293420	2+2-	INS	-103	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57299680	2+2-	20	57299695	2+2-	INS	-108	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57305083	4+1-	20	57305190	0+3-	INS	-156	31	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57311819	5+4-	20	57311924	5+4-	INS	-345	21	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57311994	2+1-	20	57312023	0+2-	INS	-169	11	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57325495	2+2-	20	57325456	2+2-	INS	-113	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57331189	2+2-	20	57331246	2+2-	INS	-187	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57347681	11+0-	20	57366706	11+1-	INV	18933	99	11	COLO-829BL-IL|3:COLO-829-IL|8	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	57352984	2+2-	20	57352982	2+2-	INS	-104	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57354366	3+0-	20	57354370	1+3-	INS	-325	33	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	57358033	2+2-	20	57358012	2+2-	INS	-116	30	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57364153	3+0-	20	57364282	7+10-	INS	-89	99	7	COLO-829BL-IL|5:COLO-829-IL|2	0.28	BreakDancerMax-0.0.1r81	|q10|o20
20	57373992	2+2-	20	57373981	2+2-	INS	-100	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	57393066	7+0-	20	57393187	1+7-	DEL	157	99	6	COLO-829BL-IL|3:COLO-829-IL|3	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	57421879	3+2-	20	57421936	3+2-	INS	-91	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57450626	2+0-	20	57450752	0+2-	DEL	88	45	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57451060	2+2-	20	57451092	2+2-	INS	-217	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57454525	2+0-	20	57454653	2+4-	INS	-139	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57461223	2+3-	20	57461235	2+3-	INS	-219	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57461871	2+3-	20	57461836	2+3-	INS	-95	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57462388	2+2-	20	57462418	2+2-	INS	-232	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57465009	2+0-	20	57464999	0+2-	INS	-221	27	2	COLO-829_v2_74|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	57530625	2+3-	20	57530611	2+3-	INS	-117	33	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57553392	4+5-	20	57553504	4+5-	INS	-242	29	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	57553823	2+2-	20	57553831	2+2-	INS	-94	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57563520	2+2-	20	57563475	2+2-	INS	-100	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57566014	2+1-	20	57566072	1+2-	INS	-255	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57576747	2+0-	20	57576970	0+3-	INS	-111	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57582185	2+0-	20	57582302	0+2-	INS	-194	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57592927	3+3-	20	57592967	3+3-	INS	-229	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57603165	2+2-	20	57603135	2+2-	INS	-236	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57634180	2+2-	20	57634160	2+2-	INS	-235	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57641504	2+2-	20	57641502	2+2-	INS	-111	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57643472	28+20-	20	57643627	28+20-	INS	-97	16	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	57647219	6+2-	20	57647475	4+4-	DEL	279	76	4	COLO-829-IL|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	57647479	0+4-	20	57647475	4+0-	ITX	-122	74	4	COLO-829BL-IL|1:COLO-829-IL|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	57666957	2+2-	20	57666951	2+2-	INS	-120	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57679149	3+3-	20	57679130	3+3-	INS	-371	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57694956	22+2-	20	57695098	22+2-	INS	-246	11	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57695168	20+0-	20	57695158	16+36-	DEL	105	99	17	COLO-829BL-IL|9:COLO-829-IL|8	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	57697913	2+2-	20	57697879	2+2-	INS	-95	36	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57700821	2+2-	20	57700830	2+2-	INS	-221	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57707013	3+0-	20	57707061	0+3-	INS	-258	30	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	57724054	2+0-	20	57724091	1+2-	INS	-301	29	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57730374	2+2-	20	57730376	2+2-	INS	-105	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	57731721	3+4-	20	57731839	0+2-	INS	-155	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57741324	2+0-	20	57741418	0+2-	INS	-227	21	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57757896	2+2-	20	57757855	2+2-	INS	-390	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57762189	2+2-	20	57762171	2+2-	INS	-104	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57770552	3+3-	20	57770628	3+3-	INS	-348	14	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57780666	3+3-	20	57780729	3+3-	INS	-240	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57789249	3+3-	20	57789241	3+3-	INS	-91	44	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57797245	2+0-	20	57797234	1+3-	INS	-268	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	57842316	3+2-	20	57842363	3+2-	INS	-228	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57844194	2+2-	20	57844145	2+2-	INS	-410	29	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	57851164	2+0-	20	57851290	1+5-	INS	-212	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57878298	2+0-	20	57878437	0+2-	INS	-191	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57879716	2+2-	20	57879705	2+2-	INS	-116	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57880955	2+2-	20	57880923	2+2-	INS	-103	32	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	57891830	2+2-	20	57891808	2+2-	INS	-99	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57893562	2+2-	20	57893511	2+2-	INS	-111	42	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	57894543	3+2-	20	57894572	3+2-	INS	-119	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57905659	3+3-	20	57905749	3+3-	INS	-186	23	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57909320	2+2-	20	57909355	2+2-	INS	-93	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57927983	3+3-	20	57928015	3+3-	INS	-111	35	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57960031	4+3-	20	57960115	4+3-	INS	-180	25	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57968178	2+2-	20	57968196	2+2-	INS	-123	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	57976486	10+12-	20	57976618	0+3-	DEL	89	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	57992589	4+2-	20	57992591	4+2-	INS	-232	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	57992661	2+0-	20	57992754	0+3-	INS	-204	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58000964	2+2-	20	58000946	2+2-	INS	-107	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58016048	3+0-	20	58016051	1+2-	INS	-346	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58073430	2+1-	20	58073413	0+2-	INS	-344	21	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	58080779	2+3-	20	58080761	2+3-	INS	-107	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58080900	3+3-	20	58080882	3+3-	INS	-289	37	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	58085712	2+3-	20	58085693	2+3-	INS	-87	33	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	58093507	2+2-	20	58093516	2+2-	INS	-111	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58102241	2+2-	20	58102273	2+2-	INS	-96	23	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	58103724	2+2-	20	58103692	2+2-	INS	-108	32	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	58106821	2+2-	20	58106908	0+2-	INS	-182	15	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58156269	2+1-	20	58156359	3+5-	INS	-258	50	5	COLO-829_v2_74|4:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	58172847	3+1-	20	58172902	0+2-	INS	-198	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58188248	2+2-	20	58188220	2+2-	INS	-378	24	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	58213859	2+2-	20	58213864	2+2-	INS	-91	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	58216725	2+2-	20	58216741	2+2-	INS	-94	29	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58222784	2+2-	20	58222745	2+2-	INS	-110	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58244515	2+2-	20	58244496	2+2-	INS	-108	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58252539	2+2-	20	58252507	2+2-	INS	-102	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	58257411	3+1-	20	58257427	0+2-	INS	-288	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58282985	3+2-	20	58283016	0+2-	INS	-157	24	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58293054	2+2-	20	58293027	2+2-	INS	-110	31	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58302079	3+0-	20	58302153	1+4-	INS	-234	51	4	COLO-829_v2_74|3:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	58322990	1+4-	20	58323094	7+4-	ITX	-97	99	6	COLO-829BL-IL|3:COLO-829_v2_74|1:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	58330892	2+2-	20	58330884	2+2-	INS	-252	21	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58336221	2+2-	20	58336175	2+2-	INS	-396	28	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58344691	9+10-	20	58344816	0+2-	INS	-132	17	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58359182	3+3-	20	58359207	1+2-	INS	-238	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58360121	34+2-	20	58360424	0+32-	DEL	327	99	29	COLO-829BL-IL|8:COLO-829_v2_74|6:COLO-829-IL|15	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	58360121	3+0-	20	58360726	0+3-	DEL	343	60	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58367712	2+2-	20	58367715	2+2-	INS	-246	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58379026	3+3-	20	58379109	3+3-	INS	-174	25	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58403895	3+2-	20	58403917	3+2-	INS	-108	23	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58412032	2+3-	20	58412024	2+3-	INS	-109	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58416137	2+1-	20	58416197	1+2-	INS	-221	14	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58421781	3+2-	20	58421798	3+2-	INS	-98	25	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58426321	2+2-	20	58426262	2+2-	INS	-115	46	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	58432968	2+0-	20	58433171	0+2-	INS	-127	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58445929	2+0-	20	58445980	1+3-	INS	-216	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	58447435	20+18-	20	58447515	20+18-	INS	-93	99	17	COLO-829BL-IL|7:COLO-829-IL|10	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	58447585	3+1-	20	58447607	0+3-	INS	-264	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58452153	3+1-	20	58452353	0+3-	INS	-141	32	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58454583	2+2-	20	58454535	2+2-	INS	-110	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58466285	2+3-	20	58466282	2+3-	INS	-260	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58469490	3+1-	20	58469512	1+2-	INS	-253	44	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	58487808	2+3-	20	58487820	2+3-	INS	-107	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58491378	2+2-	20	58491371	2+2-	INS	-114	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58498126	2+2-	20	58498073	2+2-	INS	-403	31	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58508772	2+0-	20	58509420	11+18-	DEL	368	50	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	58509356	3+14-	20	58509420	11+16-	ITX	-62	99	12	COLO-829BL-IL|5:COLO-829_v2_74|1:COLO-829-IL|6	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	58509100	16+0-	20	58509420	0+16-	DEL	344	99	16	COLO-829BL-IL|6:COLO-829-IL|10	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	58521973	2+3-	20	58521966	2+3-	INS	-105	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58526618	2+2-	20	58526647	2+2-	INS	-239	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58554537	2+2-	20	58554571	2+2-	INS	-358	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58562970	2+2-	20	58562934	2+2-	INS	-106	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58571483	4+2-	20	58571515	4+2-	INS	-102	27	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58571585	2+0-	20	58571610	0+3-	INS	-277	12	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58579353	6+4-	20	58579471	6+4-	INS	-189	23	3	COLO-829_v2_74|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58579605	2+3-	20	58579590	2+3-	INS	-108	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58588344	4+3-	20	58588405	0+3-	INS	-175	26	4	COLO-829BL-IL|1:COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58590493	3+3-	20	58590495	3+3-	INS	-115	40	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58594338	2+2-	20	58594395	2+2-	INS	-88	22	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58600859	2+1-	20	58600961	3+4-	INS	-147	34	4	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	58608651	7+6-	20	58608680	7+6-	INS	-94	87	6	COLO-829BL-IL|4:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	58617703	2+2-	20	58617695	2+2-	INS	-93	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58619672	2+2-	20	58619699	2+2-	INS	-103	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58631326	2+2-	20	58631309	2+2-	INS	-254	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58631550	2+2-	20	58631539	2+2-	INS	-227	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58636805	3+2-	20	58636867	3+2-	INS	-105	20	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58637226	3+4-	20	58637244	3+4-	INS	-118	25	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58639319	3+0-	20	58639489	0+3-	INS	-157	36	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58640351	2+2-	20	58640357	2+2-	INS	-98	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58646663	2+0-	20	58646772	1+3-	INS	-190	39	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58649638	2+2-	20	58649636	2+2-	INS	-236	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58654859	2+2-	20	58654831	2+2-	INS	-110	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58664013	2+2-	20	58664007	2+2-	INS	-248	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58674547	3+2-	20	58674536	3+2-	INS	-396	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58679384	2+0-	20	58679563	0+2-	INS	-126	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58684670	3+3-	20	58684775	3+3-	INS	-223	20	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58734192	2+3-	20	58734169	2+3-	INS	-102	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	58736944	2+2-	20	58736980	2+2-	INS	-88	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58739419	3+2-	20	58739445	3+2-	INS	-217	17	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58749395	2+2-	20	58749397	2+2-	INS	-225	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	58750929	3+4-	20	58750966	3+4-	INS	-390	27	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58764379	2+2-	20	58764360	2+2-	INS	-95	33	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58765584	2+2-	20	58765587	2+2-	INS	-100	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58768154	2+2-	20	58768123	2+2-	INS	-121	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58769042	2+0-	20	58769047	0+2-	INS	-205	29	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	58772584	73+73-	20	58773015	73+73-	DEL	89	99	56	COLO-829BL-IL|19:COLO-829-IL|37	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	58773085	3+3-	20	58773077	0+2-	DEL	78	35	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	58780683	2+3-	20	58780762	2+3-	INS	-308	13	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58782389	2+2-	20	58782402	2+2-	INS	-109	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58782607	2+2-	20	58782575	2+2-	INS	-89	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58784037	2+2-	20	58784063	2+2-	INS	-98	24	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	58785160	2+2-	20	58785191	2+2-	INS	-239	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58786818	2+1-	20	58787023	0+2-	INS	-106	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58798211	2+2-	20	58798179	2+2-	INS	-106	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58800586	7+8-	20	58800629	7+8-	INS	-91	99	7	COLO-829-IL|7	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	58803353	2+2-	20	58803394	2+2-	INS	-235	18	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58807591	3+1-	20	58807573	0+2-	INS	-217	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	58809728	2+2-	20	58809732	2+2-	INS	-106	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58840111	2+2-	20	58840106	2+2-	INS	-355	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58866791	2+2-	20	58866781	2+2-	INS	-113	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	58885312	2+2-	20	58885314	2+2-	INS	-218	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58890627	2+2-	20	58890636	2+2-	INS	-100	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58892407	3+4-	20	58892416	3+4-	INS	-257	32	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58897028	2+2-	20	58896993	2+2-	INS	-384	25	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58911507	9+11-	20	58911688	9+11-	INS	-88	48	5	COLO-829BL-IL|1:COLO-829-IL|4	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	58911758	2+4-	20	58911830	0+2-	INS	-136	9	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58919579	2+2-	20	58919555	2+2-	INS	-99	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58930289	2+2-	20	58930301	2+2-	INS	-227	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58932992	2+0-	20	58933114	0+2-	INS	-201	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	58948409	3+0-	20	58948421	0+3-	INS	-266	23	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	58956251	2+1-	20	58956272	0+2-	INS	-328	22	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	58985006	3+3-	20	58985059	3+3-	INS	-107	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59003320	5+4-	20	59003375	5+4-	INS	-363	37	4	COLO-829_v2_74|4	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	59029698	2+2-	20	59029687	2+2-	INS	-102	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59030022	2+3-	20	59030066	2+3-	INS	-103	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59031749	2+0-	20	59031920	1+4-	INS	-135	31	3	COLO-829_v2_74|2:COLO-829-IL|1	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	59034226	2+2-	20	59034196	2+2-	INS	-268	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59059985	28+0-	20	59060186	26+32-	DEL	198	99	28	COLO-829BL-IL|11:COLO-829-IL|17	0.27	BreakDancerMax-0.0.1r81	|q10|o20
20	59060204	2+25-	20	59060186	23+1-	ITX	-176	99	25	COLO-829BL-IL|9:COLO-829-IL|16	0.22	BreakDancerMax-0.0.1r81	|q10|o20
20	59068034	6+3-	20	59068142	6+3-	INS	-100	31	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59092959	3+2-	20	59093125	0+2-	INS	-128	24	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59094276	3+2-	20	59094284	3+2-	INS	-247	21	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59109431	12+0-	20	59109836	0+3-	DEL	149	45	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	59109431	10+0-	20	59109947	10+9-	DEL	233	99	9	COLO-829_v2_74|9	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	59110182	10+0-	20	59110255	44+48-	DEL	102	99	10	COLO-829BL-IL|3:COLO-829_v2_74|4:COLO-829-IL|3	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	59110747	35+30-	20	59110748	31+37-	DEL	457	99	32	COLO-829BL-IL|8:COLO-829_v2_74|4:COLO-829-IL|20	0.16	BreakDancerMax-0.0.1r81	|q10|o20
20	59110747	2+0-	20	59111272	0+2-	DEL	519	36	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59117942	2+2-	20	59117921	2+2-	INS	-257	23	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59118466	2+0-	20	59118578	0+2-	INS	-210	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59124739	4+3-	20	59124837	4+3-	INS	-255	21	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59179366	2+0-	20	59179442	0+2-	INS	-249	22	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	59181983	2+2-	20	59181986	2+2-	INS	-94	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59195443	2+2-	20	59195494	2+2-	INS	-88	21	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59196029	4+2-	20	59196046	1+3-	INS	-146	45	5	COLO-829BL-IL|2:COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	59205986	2+0-	20	59206111	1+2-	INS	-165	15	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59206091	2+2-	20	59206038	2+2-	INS	-111	37	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	59210116	3+0-	20	59210573	30+30-	ITX	-154	99	15	COLO-829BL-IL|7:COLO-829-IL|8	0.16	BreakDancerMax-0.0.1r81	|q10|o20
20	59210335	10+0-	20	59210573	14+11-	DEL	283	99	10	COLO-829BL-IL|4:COLO-829-IL|6	0.36	BreakDancerMax-0.0.1r81	|q10|o20
20	59210758	14+1-	20	59210830	0+15-	DEL	119	99	7	COLO-829BL-IL|2:COLO-829-IL|5	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	59210497	4+2-	20	59210573	2+1-	ITX	-90	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	59210497	3+0-	20	59210830	0+3-	DEL	320	54	3	COLO-829BL-IL|2:COLO-829-IL|1	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	59217375	2+2-	20	59217402	2+2-	INS	-99	28	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	59238111	2+0-	20	59238232	1+2-	DEL	89	40	2	COLO-829-IL|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	59251519	3+0-	20	59251653	0+3-	DEL	93	75	3	COLO-829BL-IL|2:COLO-829-IL|1	0.75	BreakDancerMax-0.0.1r81	|q10|o20
20	59251588	2+0-	20	59251723	0+2-	DEL	91	43	2	COLO-829-IL|2	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	59264591	3+0-	20	59264735	0+3-	INS	-172	32	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59272942	3+0-	20	59273030	19+13-	DEL	90	65	3	COLO-829BL-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59273162	19+10-	20	59273661	1+18-	DEL	519	99	18	COLO-829BL-IL|6:COLO-829-IL|12	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	59273162	1+10-	20	59273467	10+2-	ITX	135	99	10	COLO-829BL-IL|5:COLO-829-IL|5	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	59281639	17+5-	20	59281981	0+43-	DEL	265	32	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	59281639	14+4-	20	59282897	38+21-	DEL	1257	99	14	COLO-829BL-IL|6:COLO-829-IL|8	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	59281639	0+4-	20	59281757	13+4-	ITX	-17	66	4	COLO-829BL-IL|2:COLO-829-IL|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	59282252	0+41-	20	59282897	38+7-	ITX	647	99	37	COLO-829BL-IL|13:COLO-829-IL|24	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	59281998	7+2-	20	59281981	0+4-	INS	-165	20	4	COLO-829_v2_74|4	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	59281998	3+2-	20	59282897	1+7-	DEL	957	44	3	COLO-829BL-IL|2:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	59291339	12+12-	20	59291358	12+12-	INS	-101	99	10	COLO-829BL-IL|5:COLO-829-IL|5	0.16	BreakDancerMax-0.0.1r81	|q10|o20
20	59291668	7+0-	20	59291784	38+40-	INS	-151	99	17	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|13	0.27	BreakDancerMax-0.0.1r81	|q10|o20
20	59291989	8+3-	20	59292001	0+7-	INS	-176	59	7	COLO-829_v2_74|7	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	59297431	2+2-	20	59297398	2+2-	INS	-105	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59317810	2+0-	20	59317934	0+2-	DEL	93	43	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59323740	2+2-	20	59323693	2+2-	INS	-396	29	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	59334560	2+0-	20	59334749	0+2-	INS	-133	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59335462	3+2-	20	59335500	0+2-	INS	-183	26	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59337577	4+1-	20	59337567	378+381-	INS	-157	99	283	COLO-829BL-IL|76:COLO-829_v2_74|73:COLO-829-IL|134	0.74	BreakDancerMax-0.0.1r81	|q10|o20
20	59345728	10+9-	20	59345830	10+9-	INS	-227	84	9	COLO-829BL-IL|1:COLO-829_v2_74|6:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59347928	3+1-	20	59348000	1+3-	INS	-209	37	4	COLO-829_v2_74|3:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59358599	5+0-	20	59359015	0+7-	DEL	154	99	4	COLO-829_v2_74|4	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	59358813	2+1-	20	59359015	0+3-	DEL	163	38	2	COLO-829BL-IL|1:COLO-829-IL|1	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	59366497	2+0-	20	59366696	0+2-	INS	-118	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59383596	2+2-	20	59383563	2+2-	INS	-261	25	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59384031	1+2-	20	59384067	3+0-	ITX	-369	68	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	59384303	11+4-	20	59384323	11+4-	INS	-351	17	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59384393	9+2-	20	59384420	1+8-	DEL	91	99	8	COLO-829BL-IL|4:COLO-829-IL|4	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	59405944	2+0-	20	59406092	0+2-	INS	-155	20	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59437819	3+3-	20	59437898	3+3-	INS	-278	22	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59446694	2+2-	20	59446664	2+2-	INS	-93	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59452722	40+0-	20	59452719	0+40-	DEL	90	99	38	COLO-829BL-IL|17:COLO-829-IL|21	0.16	BreakDancerMax-0.0.1r81	|q10|o20
20	59454155	2+2-	20	59454141	2+2-	INS	-110	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59466368	7+20-	20	59466351	27+13-	ITX	-73	99	23	COLO-829BL-IL|2:COLO-829_v2_74|17:COLO-829-IL|4	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	59469795	2+2-	20	59469789	2+2-	INS	-89	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	59481994	2+1-	20	59482148	3+2-	INS	-194	16	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59508458	2+2-	20	59508499	2+2-	INS	-238	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	59510915	2+2-	20	59510916	2+2-	INS	-106	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59515353	2+2-	20	59515321	2+2-	INS	-381	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59526159	2+1-	20	59526163	2+3-	INS	-229	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	59527050	3+2-	20	59527153	0+3-	INS	-188	12	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59528218	3+1-	20	59528267	0+3-	INS	-195	28	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	59537843	2+2-	20	59537890	2+2-	INS	-197	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59543036	2+0-	20	59543461	0+2-	DEL	95	57	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	59543261	9+2-	20	59543271	0+9-	DEL	96	99	8	COLO-829-IL|8	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	59545209	2+2-	20	59545175	2+2-	INS	-91	36	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59554240	27+28-	20	59554695	27+28-	INS	-152	99	14	COLO-829_v2_74|14	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	59573642	4+1-	20	59573671	2+5-	DEL	90	52	3	COLO-829BL-IL|1:COLO-829-IL|2	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	59576771	2+2-	20	59576715	2+2-	INS	-120	40	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	59587285	2+2-	20	59587269	2+2-	INS	-93	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59593820	4+0-	20	59594209	1+81-	DEL	123	91	4	COLO-829_v2_74|4	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	59594181	82+4-	20	59594209	1+77-	DEL	115	99	74	COLO-829BL-IL|23:COLO-829_v2_74|4:COLO-829-IL|47	0.35	BreakDancerMax-0.0.1r81	|q10|o20
20	59594181	6+2-	20	59594487	0+6-	DEL	115	99	5	COLO-829_v2_74|5	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	59599841	3+4-	20	59599952	0+2-	INS	-150	23	3	COLO-829_v2_74|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59608814	2+2-	20	59608792	2+2-	INS	-372	23	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	59616304	2+2-	20	59616392	1+3-	INS	-267	28	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	59650146	12+2-	20	59650509	0+18-	DEL	343	99	11	COLO-829BL-IL|3:COLO-829_v2_74|3:COLO-829-IL|5	0.58	BreakDancerMax-0.0.1r81	|q10|o20
20	59650411	5+0-	20	59650509	0+7-	DEL	91	92	5	COLO-829BL-IL|3:COLO-829-IL|2	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	59676359	2+0-	20	59676451	0+2-	INS	-232	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59679100	2+2-	20	59679073	2+2-	INS	-107	31	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59684429	2+2-	20	59684399	2+2-	INS	-249	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	59698106	20+18-	20	59698173	20+18-	ITX	-170	99	16	COLO-829BL-IL|5:COLO-829-IL|11	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	59698243	4+2-	20	59698355	0+4-	INS	-177	30	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59724143	2+0-	20	59724307	0+4-	INS	-123	16	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	59752953	50+3-	20	59753259	0+2-	INS	-100	10	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59752953	46+1-	20	59752945	1+47-	DEL	125	99	46	COLO-829BL-IL|12:COLO-829_v2_74|10:COLO-829-IL|24	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	59785994	4+0-	20	59785985	42+48-	INS	-140	99	42	COLO-829BL-IL|9:COLO-829_v2_74|26:COLO-829-IL|7	0.36	BreakDancerMax-0.0.1r81	|q10|o20
20	59790853	2+3-	20	59790898	2+3-	INS	-228	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59791953	12+0-	20	59792762	1+9-	DEL	794	99	8	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|6	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	59791953	4+0-	20	59792943	1+6-	DEL	955	75	4	COLO-829BL-IL|1:COLO-829-IL|3	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	59793227	3+4-	20	59793184	3+4-	ITX	-135	77	3	COLO-829BL-IL|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59803528	23+28-	20	59803721	23+28-	INS	-189	99	22	COLO-829BL-IL|5:COLO-829_v2_74|10:COLO-829-IL|7	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	59807182	2+0-	20	59807232	0+2-	INS	-259	18	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	59814279	3+2-	20	59814319	3+2-	INS	-115	23	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59815198	2+3-	20	59815191	2+3-	INS	-116	28	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	59830781	3+3-	20	59830806	3+3-	INS	-373	17	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59831647	20+13-	20	59831899	20+13-	INS	-96	42	5	COLO-829BL-IL|2:COLO-829-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59841870	2+2-	20	59841886	2+2-	INS	-101	29	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59852779	2+2-	20	59852717	2+2-	INS	-411	37	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	59854406	2+0-	20	59854530	0+2-	INS	-205	24	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	59866779	6+2-	20	59866825	0+6-	DEL	90	99	5	COLO-829-IL|5	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59876380	2+3-	20	59876423	2+3-	INS	-247	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59886785	2+2-	20	59886804	2+2-	INS	-330	18	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	59897805	4+0-	20	59898211	24+27-	DEL	83	43	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59898414	23+24-	20	59898689	0+20-	DEL	340	99	19	COLO-829BL-IL|12:COLO-829-IL|7	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	59898414	4+24-	20	59899061	1+4-	DEL	358	70	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	59898414	1+24-	20	59898452	22+0-	ITX	-52	99	22	COLO-829BL-IL|8:COLO-829-IL|14	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	59901610	4+0-	20	59901742	0+9-	DEL	91	81	4	COLO-829-IL|4	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	59901682	4+0-	20	59901742	0+5-	DEL	90	77	4	COLO-829BL-IL|2:COLO-829-IL|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	59919537	2+4-	20	59919621	2+4-	INS	-86	24	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	59928204	56+57-	20	59928760	56+57-	INS	-302	99	30	COLO-829_v2_74|30	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	59929148	5+4-	20	59929152	5+4-	INS	-382	46	4	COLO-829_v2_74|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	59954215	5+1-	20	59956811	2+6-	DEL	2627	53	3	COLO-829BL-IL|1:COLO-829-IL|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	59955333	6+4-	20	59956811	2+3-	DEL	1465	34	2	COLO-829-IL|2	0.29	BreakDancerMax-0.0.1r81	|q10|o20
20	59955333	4+4-	20	59956953	8+4-	DEL	1733	51	3	COLO-829-IL|3	0.38	BreakDancerMax-0.0.1r81	|q10|o20
20	59955333	1+4-	20	59956590	4+9-	ITX	1123	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.29	BreakDancerMax-0.0.1r81	|q10|o20
20	59956794	2+9-	20	59956953	8+1-	ITX	60	99	8	COLO-829BL-IL|1:COLO-829-IL|7	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	59959696	5+0-	20	59960002	0+6-	DEL	297	99	5	COLO-829BL-IL|2:COLO-829-IL|3	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	59971625	3+3-	20	59971650	3+3-	INS	-276	27	3	COLO-829_v2_74|2:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	59979321	2+0-	20	59979352	16+3-	DEL	88	34	2	COLO-829-IL|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	59979550	16+1-	20	59979703	8+13-	DEL	231	99	13	COLO-829BL-IL|4:COLO-829-IL|9	0.32	BreakDancerMax-0.0.1r81	|q10|o20
20	59979550	3+1-	20	59980117	2+13-	DEL	501	52	3	COLO-829_v2_74|2:COLO-829-IL|1	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	59979919	8+0-	20	59980117	1+9-	DEL	194	99	8	COLO-829BL-IL|4:COLO-829_v2_74|1:COLO-829-IL|3	0.21	BreakDancerMax-0.0.1r81	|q10|o20
20	59986511	2+3-	20	59986516	2+3-	INS	-93	26	2	COLO-829-IL|2	0.20	BreakDancerMax-0.0.1r81	|q10|o20
20	59986955	3+2-	20	59986962	3+2-	INS	-101	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	59990306	6+5-	20	59990295	87+87-	INS	-151	99	47	COLO-829BL-IL|13:COLO-829_v2_74|14:COLO-829-IL|20	0.55	BreakDancerMax-0.0.1r81	|q10|o20
20	59993120	13+9-	20	59993233	0+4-	INS	-113	99	9	COLO-829BL-IL|2:COLO-829_v2_74|2:COLO-829-IL|5	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	60003836	3+0-	20	60004332	0+40-	DEL	309	69	3	COLO-829_v2_74|3	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	60004034	40+1-	20	60004332	0+37-	DEL	324	99	35	COLO-829BL-IL|13:COLO-829-IL|22	0.56	BreakDancerMax-0.0.1r81	|q10|o20
20	60004034	4+0-	20	60004636	0+2-	DEL	324	47	2	COLO-829_v2_74|2	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	60014250	2+0-	20	60014428	0+2-	INS	-146	22	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60027976	2+2-	20	60027964	2+2-	INS	-102	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60043562	2+7-	20	60043580	2+7-	INS	-402	18	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60054644	2+2-	20	60054603	2+2-	INS	-106	34	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60062088	2+2-	20	60062060	2+2-	INS	-99	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60067507	2+2-	20	60067504	2+2-	INS	-252	20	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	60071120	2+2-	20	60071073	2+2-	INS	-397	29	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	60077969	2+2-	20	60077915	2+2-	INS	-403	32	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60078186	2+2-	20	60078174	2+2-	INS	-381	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60091081	3+2-	20	60091080	3+2-	INS	-95	27	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60102680	2+2-	20	60102651	2+2-	INS	-102	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60106712	2+3-	20	60106774	2+3-	INS	-239	17	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60114192	22+34-	20	60114499	22+34-	INS	-137	88	12	COLO-829BL-IL|1:COLO-829_v2_74|6:COLO-829-IL|5	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	60115022	2+2-	20	60115010	2+2-	INS	-109	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60139180	2+2-	20	60139200	2+2-	INS	-234	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60142749	2+0-	20	60142804	0+2-	INS	-265	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60147911	2+2-	20	60147953	2+2-	INS	-239	16	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60173749	2+2-	20	60173744	2+2-	INS	-105	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60216041	2+2-	20	60216047	2+2-	INS	-97	26	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60234881	2+3-	20	60234847	2+3-	INS	-109	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60249069	2+2-	20	60249082	2+2-	INS	-219	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60263347	3+0-	20	60263444	0+2-	INS	-207	19	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60278888	7+1-	20	60278933	1+4-	DEL	87	66	4	COLO-829BL-IL|1:COLO-829-IL|3	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	60278888	2+0-	20	60279408	0+4-	DEL	250	45	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	60286661	12+0-	20	60287139	11+50-	DEL	641	99	11	COLO-829BL-IL|7:COLO-829-IL|4	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	60287105	45+8-	20	60287139	9+37-	DEL	144	99	35	COLO-829BL-IL|14:COLO-829_v2_74|2:COLO-829-IL|19	0.16	BreakDancerMax-0.0.1r81	|q10|o20
20	60286806	2+0-	20	60287139	1+2-	DEL	132	42	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	60287105	10+0-	20	60287442	0+11-	DEL	151	99	10	COLO-829_v2_74|10	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	60292503	2+2-	20	60292486	2+2-	INS	-97	33	2	COLO-829BL-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60347311	2+2-	20	60347295	2+2-	INS	-251	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	60361083	2+2-	20	60361055	2+2-	INS	-245	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60381922	3+2-	20	60382331	0+2-	DEL	140	47	2	COLO-829_v2_74|2	0.40	BreakDancerMax-0.0.1r81	|q10|o20
20	60390715	7+9-	20	60390755	7+9-	INS	-95	64	5	COLO-829BL-IL|2:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60394859	2+2-	20	60394841	2+2-	INS	-244	22	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60415080	3+0-	20	60415207	0+3-	DEL	90	62	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60420021	2+2-	20	60419984	2+2-	INS	-98	33	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	60426274	2+2-	20	60426437	0+4-	DEL	150	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	60426274	0+2-	20	60426269	5+1-	ITX	-179	53	3	COLO-829BL-IL|1:COLO-829-IL|2	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	60434551	2+0-	20	60434685	0+2-	DEL	88	50	2	COLO-829BL-IL|1:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	60454612	3+5-	20	60454574	3+5-	INS	-108	52	3	COLO-829BL-IL|2:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	60475260	2+2-	20	60475256	2+2-	INS	-106	26	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60475674	2+2-	20	60475625	2+2-	INS	-399	29	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60490796	2+2-	20	60490754	2+2-	INS	-105	34	2	COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	60505556	2+3-	20	60505619	2+3-	INS	-228	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60507230	3+0-	20	60507365	0+3-	DEL	100	69	3	COLO-829BL-IL|1:COLO-829-IL|2	0.38	BreakDancerMax-0.0.1r81	|q10|o20
20	60512829	8+10-	20	60512968	8+10-	INS	-142	56	6	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|4	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60517669	8+0-	20	60517718	0+8-	DEL	92	99	8	COLO-829BL-IL|2:COLO-829-IL|6	0.32	BreakDancerMax-0.0.1r81	|q10|o20
20	60576627	2+2-	20	60576603	2+2-	INS	-382	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60579922	2+2-	20	60579939	2+2-	INS	-235	20	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	60581569	2+2-	20	60581518	2+2-	INS	-113	38	2	COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	60587277	24+10-	20	60587301	19+35-	ITX	-75	99	21	COLO-829BL-IL|5:COLO-829-IL|16	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	60587277	2+0-	20	60587613	0+2-	DEL	488	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60605586	2+0-	20	60605649	0+3-	INS	-227	18	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	60621434	2+2-	20	60621446	2+2-	INS	-108	25	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	60741311	3+3-	20	60741352	3+3-	INS	-98	34	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60757029	2+0-	20	60757116	0+2-	DEL	93	37	2	COLO-829BL-IL|1:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	60764880	2+2-	20	60764856	2+2-	INS	-107	30	2	COLO-829-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	60774695	17+0-	20	60775583	0+17-	DEL	894	99	17	COLO-829BL-IL|9:COLO-829-IL|8	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	60778210	2+2-	20	60778193	2+2-	INS	-243	24	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	60785827	3+0-	20	60785955	0+3-	DEL	88	70	3	COLO-829BL-IL|1:COLO-829-IL|2	0.21	BreakDancerMax-0.0.1r81	|q10|o20
20	60787627	2+2-	20	60787641	2+2-	INS	-106	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60800654	24+0-	20	60800697	0+25-	DEL	103	99	22	COLO-829BL-IL|9:COLO-829-IL|13	0.19	BreakDancerMax-0.0.1r81	|q10|o20
20	60818306	9+8-	20	60818366	9+8-	INS	-98	99	8	COLO-829BL-IL|4:COLO-829-IL|4	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	60841790	3+3-	20	60841869	3+3-	INS	-198	24	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60871025	2+2-	20	60870994	2+2-	INS	-251	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60899112	3+0-	20	60899108	0+3-	INS	-333	20	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	60923352	3+3-	20	60923333	3+3-	INS	-280	35	3	COLO-829_v2_74|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	60925951	2+0-	20	60926018	4+7-	INS	-95	29	3	COLO-829BL-IL|2:COLO-829-IL|1	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	60933561	2+0-	20	60933678	0+3-	INS	-203	20	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	60941494	34+0-	20	60941820	1+6-	DEL	102	99	5	COLO-829_v2_74|5	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	60941494	29+0-	20	60941539	0+31-	DEL	106	99	29	COLO-829BL-IL|11:COLO-829-IL|18	0.51	BreakDancerMax-0.0.1r81	|q10|o20
20	60960253	2+0-	20	60960372	3+4-	INS	-126	25	3	COLO-829_v2_74|2:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60960514	2+1-	20	60960704	0+2-	DEL	92	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60961130	2+0-	20	60961112	0+3-	INS	-322	20	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	60971185	1+3-	20	60971722	0+3-	INV	298	60	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	60988514	2+2-	20	60988472	2+2-	INS	-106	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61023200	2+3-	20	61023218	2+3-	INS	-354	18	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61023639	2+2-	20	61023628	2+2-	INS	-91	27	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61025861	2+2-	20	61025858	2+2-	INS	-232	22	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61035180	2+2-	20	61035139	2+2-	INS	-116	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61041402	2+3-	20	61041433	2+3-	INS	-97	22	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61057416	2+2-	20	61057426	2+2-	INS	-231	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61068158	2+3-	20	61068120	2+3-	INS	-115	33	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61073580	8+14-	20	61073714	19+15-	ITX	-21	99	19	COLO-829BL-IL|10:COLO-829-IL|9	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	61073580	6+2-	20	61074061	0+6-	DEL	453	99	6	COLO-829BL-IL|3:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61073580	0+2-	20	61073600	5+0-	ITX	-367	55	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61073727	3+0-	20	61073714	0+6-	INS	-166	18	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61077605	3+0-	20	61077934	0+13-	DEL	81	69	3	COLO-829_v2_74|3	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	61077892	13+0-	20	61077934	0+10-	DEL	132	99	9	COLO-829BL-IL|4:COLO-829-IL|5	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	61077892	4+0-	20	61078173	0+4-	DEL	91	68	3	COLO-829_v2_74|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	61092031	2+2-	20	61092095	0+2-	DEL	87	36	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61095472	3+0-	20	61095603	0+3-	DEL	92	75	3	COLO-829BL-IL|2:COLO-829-IL|1	0.60	BreakDancerMax-0.0.1r81	|q10|o20
20	61104936	4+4-	20	61105029	4+4-	INS	-102	24	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61106689	2+1-	20	61106671	1+3-	INS	-172	30	3	COLO-829BL-IL|2:COLO-829_v2_74|1	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	61117759	7+7-	20	61117815	7+7-	INS	-94	78	6	COLO-829BL-IL|3:COLO-829-IL|3	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	61127327	2+2-	20	61127319	2+2-	INS	-113	28	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61131138	4+5-	20	61131161	4+5-	INS	-106	52	4	COLO-829BL-IL|1:COLO-829-IL|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61150798	14+6-	20	61150886	14+6-	INS	-95	24	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61170390	4+3-	20	61170345	4+3-	INS	-207	46	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	61194078	3+3-	20	61194083	3+3-	INS	-88	41	3	COLO-829BL-IL|2:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61194998	4+1-	20	61196040	1+37-	INS	-92	20	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61195181	36+1-	20	61196040	0+34-	DEL	905	99	33	COLO-829BL-IL|14:COLO-829-IL|19	0.97	BreakDancerMax-0.0.1r81	|q10|o20
20	61195181	2+0-	20	61196377	0+2-	DEL	915	46	2	COLO-829_v2_74|2	0.67	BreakDancerMax-0.0.1r81	|q10|o20
20	61203444	7+13-	20	61203666	7+13-	DEL	91	65	4	COLO-829-IL|4	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	61210670	2+3-	20	61210685	2+3-	INS	-107	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	61217838	3+3-	20	61217819	3+3-	INS	-211	39	3	COLO-829_v2_74|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61231390	2+0-	20	61231421	0+2-	INS	-288	21	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61236451	4+0-	20	61236961	0+5-	DEL	470	98	4	COLO-829BL-IL|3:COLO-829-IL|1	0.67	BreakDancerMax-0.0.1r81	|q10|o20
20	61238192	2+0-	20	61238178	0+2-	INS	-322	18	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	61240333	2+0-	20	61240343	0+3-	INS	-307	19	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61245089	2+2-	20	61245047	2+2-	INS	-113	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61248507	2+3-	20	61248576	2+3-	INS	-195	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61258657	17+0-	20	61258944	7+26-	DEL	144	99	17	COLO-829_v2_74|17	0.49	BreakDancerMax-0.0.1r81	|q10|o20
20	61258821	2+0-	20	61258944	0+2-	DEL	90	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	61272860	2+0-	20	61272982	1+2-	INS	-182	22	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61291422	2+0-	20	61291411	3+5-	INS	-162	45	5	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	61296514	7+1-	20	61299730	9+9-	DEL	3250	99	7	COLO-829BL-IL|2:COLO-829-IL|5	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	61296745	1+10-	20	61299730	9+2-	ITX	2855	99	9	COLO-829BL-IL|4:COLO-829-IL|5	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	61298130	2+2-	20	61298098	2+2-	INS	-108	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	61308586	6+3-	20	61308607	2+4-	INS	-268	52	7	COLO-829_v2_74|5:COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61320908	2+2-	20	61320878	2+2-	INS	-244	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61322595	3+2-	20	61322556	3+2-	INS	-124	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61323400	20+0-	20	61323714	1+3-	DEL	133	67	3	COLO-829_v2_74|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	61323400	17+0-	20	61323436	1+20-	DEL	115	99	17	COLO-829BL-IL|6:COLO-829-IL|11	0.26	BreakDancerMax-0.0.1r81	|q10|o20
20	61340699	2+3-	20	61340679	2+3-	INS	-101	29	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61368648	3+0-	20	61368723	0+3-	DEL	90	53	3	COLO-829BL-IL|1:COLO-829-IL|2	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	61405892	27+27-	20	61406035	27+27-	INS	-109	99	17	COLO-829BL-IL|9:COLO-829-IL|8	0.27	BreakDancerMax-0.0.1r81	|q10|o20
20	61415217	2+2-	20	61415186	2+2-	INS	-87	30	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61433994	2+3-	20	61434019	2+3-	INS	-107	24	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61458963	3+0-	20	61459059	0+3-	DEL	94	57	3	COLO-829BL-IL|1:COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	61474025	3+1-	20	61474326	3+5-	INS	-93	48	4	COLO-829BL-IL|2:COLO-829-IL|2	0.17	BreakDancerMax-0.0.1r81	|q10|o20
20	61494157	2+0-	20	61494542	0+10-	DEL	90	47	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61494486	8+0-	20	61494542	0+8-	DEL	94	99	8	COLO-829BL-IL|3:COLO-829-IL|5	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	61505311	3+2-	20	61505321	3+2-	INS	-235	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61517678	3+0-	20	61517709	0+3-	INS	-281	35	3	COLO-829_v2_74|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	61531026	2+2-	20	61531042	2+2-	INS	-242	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61533897	4+5-	20	61533866	4+5-	INS	-109	67	4	COLO-829BL-IL|1:COLO-829-IL|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	61534517	15+5-	20	61534637	0+10-	DEL	120	99	10	COLO-829BL-IL|3:COLO-829-IL|7	0.19	BreakDancerMax-0.0.1r81	|q10|o20
20	61539010	2+0-	20	61539174	0+2-	INS	-172	27	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61544576	8+1-	20	61544663	14+9-	DEL	87	70	5	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|3	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	61544681	7+1-	20	61545037	15+14-	INS	-170	23	4	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	61547679	2+1-	20	61547742	2+3-	DEL	88	35	2	COLO-829BL-IL|1:COLO-829-IL|1	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	61557578	7+0-	20	61557676	2+7-	DEL	101	99	7	COLO-829BL-IL|1:COLO-829-IL|6	0.30	BreakDancerMax-0.0.1r81	|q10|o20
20	61557834	2+0-	20	61557936	0+2-	DEL	87	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	61569152	4+4-	20	61569153	4+4-	INS	-97	57	4	COLO-829BL-IL|2:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61577651	2+2-	20	61577675	2+2-	INS	-235	19	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61581273	2+2-	20	61581299	2+2-	INS	-354	17	2	COLO-829_v2_74|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	61588780	23+22-	20	61588910	8+9-	INS	-114	99	15	COLO-829BL-IL|4:COLO-829_v2_74|1:COLO-829-IL|10	0.19	BreakDancerMax-0.0.1r81	|q10|o20
20	61588780	0+2-	20	61588771	2+2-	ITX	-179	31	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61588919	0+2-	20	61588910	2+0-	ITX	-186	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	61593919	4+6-	20	61593907	46+48-	ITX	-171	99	17	COLO-829BL-IL|3:COLO-829_v2_74|6:COLO-829-IL|8	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	61594429	11+9-	20	61594534	0+4-	DEL	260	37	3	COLO-829BL-IL|1:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61594429	8+9-	20	61594418	5+7-	DEL	90	91	6	COLO-829-IL|6	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61635495	2+3-	20	61635466	2+3-	INS	-258	24	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	61645527	2+2-	20	61645491	2+2-	INS	-102	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61661280	8+1-	20	61661578	0+8-	DEL	288	99	7	COLO-829BL-IL|1:COLO-829-IL|6	0.50	BreakDancerMax-0.0.1r81	|q10|o20
20	61663798	2+2-	20	61663763	2+2-	INS	-104	32	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61668266	65+65-	20	61668527	65+65-	INS	-143	99	41	COLO-829BL-IL|9:COLO-829_v2_74|7:COLO-829-IL|25	0.21	BreakDancerMax-0.0.1r81	|q10|o20
20	61672984	5+0-	20	61673023	12+10-	DEL	105	38	2	COLO-829BL-IL|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	61673163	10+6-	20	61673196	27+17-	DEL	90	65	4	COLO-829BL-IL|1:COLO-829-IL|3	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	61673163	6+5-	20	61673727	24+43-	INS	-247	46	6	COLO-829BL-IL|1:COLO-829_v2_74|3:COLO-829-IL|2	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	61673163	2+5-	20	61673520	9+4-	ITX	193	97	5	COLO-829BL-IL|2:COLO-829_v2_74|1:COLO-829-IL|2	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	61673425	26+13-	20	61673727	16+31-	DEL	398	99	26	COLO-829BL-IL|10:COLO-829-IL|16	0.70	BreakDancerMax-0.0.1r81	|q10|o20
20	61673933	5+5-	20	61673932	0+4-	INS	-200	27	4	COLO-829_v2_74|4	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	61673688	4+2-	20	61673727	1+5-	INS	-192	10	2	COLO-829_v2_74|2	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	61681866	4+0-	20	61682059	3+5-	DEL	163	92	4	COLO-829BL-IL|2:COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61352956	11+0-	20	61716517	7+4-	INV	363497	99	7	COLO-829-IL|7	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	61682149	2+0-	20	61682323	0+2-	INS	-164	24	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61690907	2+2-	20	61690891	2+2-	INS	-106	33	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	61708966	10+1-	20	61711272	37+64-	DEL	1155	99	18	COLO-829BL-IL|10:COLO-829-IL|8	0.23	BreakDancerMax-0.0.1r81	|q10|o20
20	61708966	2+1-	20	61708993	29+14-	DEL	88	31	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61711287	15+7-	20	61711272	26+45-	DEL	138	35	3	COLO-829BL-IL|1:COLO-829-IL|2	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	61709166	28+11-	20	61711272	26+42-	DEL	2199	99	13	COLO-829BL-IL|2:COLO-829-IL|11	0.30	BreakDancerMax-0.0.1r81	|q10|o20
20	61711082	9+9-	20	61711272	21+29-	ITX	166	38	3	COLO-829BL-IL|1:COLO-829-IL|2	0.19	BreakDancerMax-0.0.1r81	|q10|o20
20	61710699	33+44-	20	61711272	18+29-	ITX	232	99	13	COLO-829BL-IL|5:COLO-829-IL|8	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	61710990	74+82-	20	61711272	11+22-	ITX	-46	99	23	COLO-829BL-IL|9:COLO-829_v2_74|3:COLO-829-IL|11	0.27	BreakDancerMax-0.0.1r81	|q10|o20
20	61709476	37+24-	20	61711272	5+5-	ITX	1477	90	6	COLO-829-IL|6	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	61709166	14+5-	20	61710556	18+29-	ITX	1296	70	4	COLO-829BL-IL|1:COLO-829-IL|3	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	61709166	10+1-	20	61710764	29+48-	DEL	1647	99	8	COLO-829BL-IL|2:COLO-829-IL|6	0.21	BreakDancerMax-0.0.1r81	|q10|o20
20	61710990	29+40-	20	61711108	10+5-	DEL	176	81	5	COLO-829BL-IL|1:COLO-829-IL|4	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	61710699	14+25-	20	61711108	8+0-	ITX	254	99	7	COLO-829BL-IL|3:COLO-829-IL|4	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	61709476	32+18-	20	61711000	8+5-	ITX	1373	84	4	COLO-829BL-IL|1:COLO-829-IL|3	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	61710699	14+18-	20	61711000	4+1-	ITX	118	45	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61710276	4+3-	20	61710556	14+16-	ITX	162	57	3	COLO-829BL-IL|1:COLO-829-IL|2	0.33	BreakDancerMax-0.0.1r81	|q10|o20
20	61710699	11+15-	20	61710764	24+38-	ITX	-49	99	10	COLO-829BL-IL|3:COLO-829-IL|7	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	61709476	28+14-	20	61710556	1+5-	DEL	1120	73	4	COLO-829BL-IL|1:COLO-829-IL|3	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	61710276	3+0-	20	61710764	14+28-	DEL	450	51	3	COLO-829BL-IL|2:COLO-829-IL|1	0.33	BreakDancerMax-0.0.1r81	|q10|o20
20	61709476	24+13-	20	61710764	14+25-	DEL	1328	99	24	COLO-829BL-IL|12:COLO-829-IL|12	0.40	BreakDancerMax-0.0.1r81	|q10|o20
20	61709648	2+2-	20	61709765	0+2-	DEL	90	40	2	COLO-829BL-IL|1:COLO-829-IL|1	0.40	BreakDancerMax-0.0.1r81	|q10|o20
20	61715141	2+2-	20	61715087	2+2-	INS	-119	39	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61719528	13+11-	20	61719571	0+2-	INS	-116	99	12	COLO-829BL-IL|1:COLO-829_v2_74|2:COLO-829-IL|9	0.16	BreakDancerMax-0.0.1r81	|q10|o20
20	61720915	2+2-	20	61720918	2+2-	INS	-93	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61733961	0+2-	20	61740623	4+5-	INV	6543	58	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	61757695	2+3-	20	61757655	2+3-	INS	-107	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61780677	2+2-	20	61780658	2+2-	INS	-114	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61790893	2+2-	20	61790894	2+2-	INS	-108	27	2	COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	61824318	4+5-	20	61824432	4+5-	INS	-195	22	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61825334	3+0-	20	61825469	0+3-	DEL	89	75	3	COLO-829-IL|3	0.43	BreakDancerMax-0.0.1r81	|q10|o20
20	61833320	109+2-	20	61833568	2+23-	DEL	113	99	21	COLO-829_v2_74|21	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	61833320	87+1-	20	61833355	1+87-	DEL	101	99	87	COLO-829BL-IL|38:COLO-829_v2_74|7:COLO-829-IL|42	0.23	BreakDancerMax-0.0.1r81	|q10|o20
20	61834092	2+4-	20	61834145	2+4-	INS	-249	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	61859675	19+2-	20	61859736	4+21-	DEL	117	99	18	COLO-829BL-IL|6:COLO-829-IL|12	0.26	BreakDancerMax-0.0.1r81	|q10|o20
20	61864837	4+4-	20	61864880	4+4-	INS	-113	36	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61871568	2+2-	20	61871574	2+2-	INS	-95	30	2	COLO-829BL-IL|2	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	61872443	3+0-	20	61872823	0+17-	DEL	95	70	3	COLO-829_v2_74|3	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	61872784	16+0-	20	61872823	0+14-	DEL	92	99	12	COLO-829BL-IL|6:COLO-829-IL|6	0.19	BreakDancerMax-0.0.1r81	|q10|o20
20	61872784	3+0-	20	61873069	1+2-	DEL	84	45	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	61817911	0+2-	20	61908986	2+0-	ITX	90897	42	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	61933643	2+2-	20	61933605	2+2-	INS	-108	33	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61937490	2+0-	20	61937528	1+3-	INS	-209	25	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	61944339	3+3-	20	61944386	3+3-	INS	-269	27	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61948843	65+66-	20	61949367	65+66-	INS	-110	99	57	COLO-829BL-IL|17:COLO-829_v2_74|21:COLO-829-IL|19	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	61951672	20+3-	20	61951953	6+2-	DEL	92	43	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	61951672	18+3-	20	61951725	0+18-	DEL	102	99	18	COLO-829BL-IL|4:COLO-829-IL|14	0.30	BreakDancerMax-0.0.1r81	|q10|o20
20	61970960	3+2-	20	61970944	3+2-	INS	-106	29	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61994631	5+2-	20	61994687	5+2-	INS	-202	15	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	61999725	3+3-	20	61999760	3+3-	INS	-386	16	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62000995	3+3-	20	62001065	3+3-	INS	-374	24	3	COLO-829_v2_74|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62010465	2+2-	20	62010440	2+2-	INS	-375	23	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62014967	24+19-	20	62015078	2+4-	INS	-169	99	20	COLO-829BL-IL|5:COLO-829_v2_74|6:COLO-829-IL|9	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	62021670	2+0-	20	62022082	0+2-	DEL	79	58	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62050418	2+2-	20	62050436	2+2-	INS	-230	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	62066653	26+0-	20	62068201	0+3-	DEL	1267	75	3	COLO-829_v2_74|3	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	62066653	23+0-	20	62067917	0+24-	DEL	1281	99	23	COLO-829BL-IL|8:COLO-829-IL|15	0.26	BreakDancerMax-0.0.1r81	|q10|o20
20	62072744	43+32-	20	62072733	0+14-	INS	-141	99	35	COLO-829BL-IL|7:COLO-829_v2_74|14:COLO-829-IL|14	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	62087187	2+0-	20	62087277	0+2-	INS	-232	21	2	COLO-829_v2_74|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62090423	3+2-	20	62090458	3+2-	INS	-92	23	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62128664	3+2-	20	62128628	3+2-	INS	-111	33	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62136646	2+2-	20	62136663	2+2-	INS	-240	18	2	COLO-829_v2_74|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62161837	3+1-	20	62161990	0+2-	INS	-127	31	3	COLO-829BL-IL|1:COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62179993	22+21-	20	62180042	22+21-	INS	-95	99	20	COLO-829BL-IL|5:COLO-829-IL|15	0.12	BreakDancerMax-0.0.1r81	|q10|o20
20	62190286	5+1-	20	62190274	128+133-	INS	-122	99	51	COLO-829BL-IL|11:COLO-829_v2_74|5:COLO-829-IL|35	0.26	BreakDancerMax-0.0.1r81	|q10|o20
20	62190539	58+60-	20	62190535	156+155-	ITX	-153	99	119	COLO-829BL-IL|30:COLO-829_v2_74|9:COLO-829-IL|80	0.26	BreakDancerMax-0.0.1r81	|q10|o20
20	62192584	4+0-	20	62193242	0+3-	DEL	321	84	3	COLO-829_v2_74|3	0.50	BreakDancerMax-0.0.1r81	|q10|o20
20	62198712	6+2-	20	62198776	11+13-	INS	-284	76	8	COLO-829_v2_74|8	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	62199200	3+3-	20	62199165	3+3-	INS	-104	31	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	62206171	2+3-	20	62206175	2+3-	INS	-102	30	2	COLO-829BL-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	62219233	2+1-	20	62220314	7+6-	ITX	383	32	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	62220276	3+3-	20	62220314	5+4-	DEL	88	48	3	COLO-829BL-IL|1:COLO-829-IL|2	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	62219644	1+6-	20	62220314	4+1-	ITX	536	33	2	COLO-829BL-IL|1:COLO-829-IL|1	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	62220033	1+2-	20	62220886	3+1-	ITX	445	62	3	COLO-829BL-IL|2:COLO-829-IL|1	0.23	BreakDancerMax-0.0.1r81	|q10|o20
20	62225050	18+20-	20	62225054	32+1-	ITX	-92	99	19	COLO-829BL-IL|9:COLO-829-IL|10	0.15	BreakDancerMax-0.0.1r81	|q10|o20
20	62225050	17+0-	20	62225289	16+45-	DEL	277	99	17	COLO-829BL-IL|2:COLO-829-IL|15	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	62225208	12+0-	20	62225289	0+12-	DEL	93	99	12	COLO-829BL-IL|5:COLO-829-IL|7	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	62227010	6+5-	20	62227167	6+5-	INS	-94	28	3	COLO-829BL-IL|2:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62227237	3+2-	20	62227533	0+2-	DEL	332	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62228039	14+1-	20	62228371	0+14-	DEL	347	99	14	COLO-829BL-IL|6:COLO-829-IL|8	0.21	BreakDancerMax-0.0.1r81	|q10|o20
20	62233096	2+2-	20	62233079	2+2-	INS	-97	28	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62233910	23+8-	20	62233909	40+40-	DEL	267	99	18	COLO-829BL-IL|5:COLO-829-IL|13	0.31	BreakDancerMax-0.0.1r81	|q10|o20
20	62233910	13+1-	20	62234785	5+9-	DEL	1084	75	5	COLO-829BL-IL|2:COLO-829-IL|3	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	62233910	8+1-	20	62234682	4+8-	DEL	1062	42	3	COLO-829BL-IL|2:COLO-829-IL|1	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	62233910	5+1-	20	62235658	0+16-	DEL	1739	55	4	COLO-829BL-IL|1:COLO-829-IL|3	0.09	BreakDancerMax-0.0.1r81	|q10|o20
20	62234590	14+11-	20	62234592	8+5-	ITX	244	27	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62234590	12+9-	20	62235478	2+2-	DEL	1002	21	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62234590	10+9-	20	62235658	0+12-	DEL	1125	35	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	62234590	7+9-	20	62234785	5+4-	ITX	212	63	5	COLO-829BL-IL|1:COLO-829-IL|4	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	62234590	4+4-	20	62234682	4+5-	DEL	255	47	4	COLO-829BL-IL|2:COLO-829-IL|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	62234690	4+1-	20	62235658	0+9-	DEL	958	65	3	COLO-829BL-IL|3	0.38	BreakDancerMax-0.0.1r81	|q10|o20
20	62235491	2+0-	20	62235658	0+6-	DEL	196	43	2	COLO-829BL-IL|2	1.00	BreakDancerMax-0.0.1r81	|q10|o20
20	62235595	2+0-	20	62235658	0+4-	DEL	90	34	2	COLO-829BL-IL|1:COLO-829-IL|1	0.10	BreakDancerMax-0.0.1r81	|q10|o20
20	62236753	2+0-	20	62237244	27+11-	DEL	183	43	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	62237512	27+9-	20	62237719	3+26-	DEL	315	99	25	COLO-829BL-IL|9:COLO-829-IL|16	0.17	BreakDancerMax-0.0.1r81	|q10|o20
20	62236864	2+0-	20	62237244	2+9-	DEL	202	42	2	COLO-829_v2_74|2	0.08	BreakDancerMax-0.0.1r81	|q10|o20
20	62236976	8+0-	20	62237244	2+7-	DEL	149	99	5	COLO-829_v2_74|4:COLO-829-IL|1	0.45	BreakDancerMax-0.0.1r81	|q10|o20
20	62237175	2+0-	20	62237244	2+2-	DEL	86	29	2	COLO-829BL-IL|1:COLO-829-IL|1	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	62237512	2+0-	20	62238052	1+2-	DEL	310	41	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62237936	3+1-	20	62238294	0+7-	DEL	82	65	3	COLO-829_v2_74|3	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62236976	3+0-	20	62237494	0+2-	DEL	209	52	2	COLO-829_v2_74|2	0.25	BreakDancerMax-0.0.1r81	|q10|o20
20	62238267	3+0-	20	62238294	0+4-	DEL	87	40	2	COLO-829BL-IL|2	0.06	BreakDancerMax-0.0.1r81	|q10|o20
20	62249314	3+4-	20	62249345	3+4-	INS	-97	45	3	COLO-829BL-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62251753	2+0-	20	62251850	2+6-	INS	-121	28	3	COLO-829BL-IL|1:COLO-829_v2_74|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	62255733	2+1-	20	62255809	0+4-	INS	-233	18	2	COLO-829_v2_74|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	62260052	6+0-	20	62260156	0+6-	DEL	103	99	6	COLO-829BL-IL|1:COLO-829-IL|5	0.23	BreakDancerMax-0.0.1r81	|q10|o20
20	62266560	2+2-	20	62266528	2+2-	INS	-96	32	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62268450	2+0-	20	62268491	0+2-	INS	-276	20	2	COLO-829_v2_74|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62270554	2+2-	20	62270557	2+2-	INS	-111	25	2	COLO-829BL-IL|1:COLO-829-IL|1	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	62275572	52+55-	20	62277697	9+1-	INS	-105	99	31	COLO-829BL-IL|10:COLO-829-IL|21	0.60	BreakDancerMax-0.0.1r81	|q10|o20
20	62275572	6+3-	20	62278026	4+14-	DEL	2566	99	6	COLO-829BL-IL|2:COLO-829-IL|4	0.22	BreakDancerMax-0.0.1r81	|q10|o20
20	62277794	2+0-	20	62277832	7+2-	DEL	85	34	2	COLO-829-IL|2	0.18	BreakDancerMax-0.0.1r81	|q10|o20
20	62278020	7+0-	20	62278026	2+6-	DEL	90	99	6	COLO-829BL-IL|2:COLO-829-IL|4	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	62280452	19+20-	20	62280451	0+2-	INS	-143	99	16	COLO-829BL-IL|6:COLO-829_v2_74|6:COLO-829-IL|4	0.11	BreakDancerMax-0.0.1r81	|q10|o20
20	62280452	0+3-	20	62280903	3+0-	ITX	330	45	3	COLO-829BL-IL|1:COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62286980	2+0-	20	62287061	0+2-	INS	-242	22	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	62299172	2+2-	20	62299248	2+2-	INS	-180	16	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62303827	5+4-	20	62303844	5+4-	ITX	-134	39	2	COLO-829-IL|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	62309992	3+2-	20	62309967	3+2-	INS	-394	23	2	COLO-829_v2_74|2	0.03	BreakDancerMax-0.0.1r81	|q10|o20
20	62314684	2+2-	20	62314694	2+2-	INS	-94	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62325496	2+2-	20	62325505	2+2-	INS	-101	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62331578	2+2-	20	62331553	2+2-	INS	-375	23	2	COLO-829_v2_74|2	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	62338411	2+2-	20	62338416	2+2-	INS	-237	19	2	COLO-829_v2_74|1:COLO-829-IL|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	62346062	2+2-	20	62346034	2+2-	INS	-246	26	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	62349879	2+2-	20	62349899	2+2-	INS	-94	29	2	COLO-829BL-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62351993	3+4-	20	62352123	3+4-	INS	-90	36	3	COLO-829BL-IL|3	0.01	BreakDancerMax-0.0.1r81	|q10|o20
20	62356919	2+3-	20	62356906	2+3-	INS	-114	28	2	COLO-829-IL|2	0.02	BreakDancerMax-0.0.1r81	|q10|o20
20	62369424	2+2-	20	62369417	2+2-	INS	-220	23	2	COLO-829BL-IL|1:COLO-829_v2_74|1	0.00	BreakDancerMax-0.0.1r81	|q10|o20
20	62372515	5+2-	20	62372516	5+2-	INS	-96	27	2	COLO-829-IL|2	0.05	BreakDancerMax-0.0.1r81	|q10|o20
20	62372586	3+0-	20	62373285	0+3-	DEL	374	78	3	COLO-829_v2_74|3	0.07	BreakDancerMax-0.0.1r81	|q10|o20
20	62388719	7+14-	20	62389050	58+138-	ITX	324	24	2	COLO-829BL-IL|1:COLO-829-IL|1	0.04	BreakDancerMax-0.0.1r81	|q10|o20
20	62388719	6+11-	20	62388756	47+52-	DEL	90	99	7	COLO-829BL-IL|2:COLO-829-IL|5	0.14	BreakDancerMax-0.0.1r81	|q10|o20
20	62389053	43+44-	20	62389050	54+136-	DEL	116	99	26	COLO-829BL-IL|9:COLO-829_v2_74|1:COLO-829-IL|16	0.13	BreakDancerMax-0.0.1r81	|q10|o20
20	62416081	2+2-	20	62416055	2+2-	INS	-126	31	2	COLO-829-IL|2	0.01	BreakDancerMax-0.0.1r81	|q10|o20
